module FIFO_in(input0, output0, output1, output2, output3, output4, output5, output6, output7, output8, output9, output10, output11, output12, output13, output14, output15, command, col, resetn,clk);
input [31:0] input0;
input [1:0] command;
input [1:0] col;
output [7:0] output0, output1, output2, output3, output4, output5, output6, output7, output8, output9, output10, output11, output12, output13, output14, output15;
input clk , resetn;

/*reg signed [23:0] x0,x1,x2,x3,x4,x5,x6,x7;
reg signed [24:0] a0,a1,a2,a3,b0,b1,b2,b3;
reg signed [30:0] m0_64,m1_64,m2_64,m3_64;
reg signed [28:0] m0_9,m1_9,m2_9,m3_9;
reg signed [29:0] m0_25,m1_25,m2_25,m3_25;
reg signed [31:0] t0_18,t0_50,t0_75,t0_89,t1_18,t1_50,t1_75,t1_89,t2_18,t2_50,t2_75,t2_89,t3_18,t3_50,t3_75,t3_89;
reg signed [32:0] stageI [0:7];
reg signed [33:0] y1,y3,y5,y7;
wire signed [23:0] y0,y2,y4,y6;*/

wire load_enable, fifo_enable;
reg [7:0]  in_reg0_0, in_reg1_0, in_reg1_1, in_reg2_0, in_reg2_1, in_reg2_2, in_reg3_0, in_reg3_1, in_reg3_2, in_reg3_3, in_reg4_0, in_reg4_1, in_reg4_2, in_reg4_3, in_reg4_4, in_reg5_0, in_reg5_1, in_reg5_2, in_reg5_3, in_reg5_4, in_reg5_5, in_reg6_0, in_reg6_1, in_reg6_2, in_reg6_3, in_reg6_4, in_reg6_5, in_reg6_6, in_reg7_0, in_reg7_1, in_reg7_2, in_reg7_3, in_reg7_4, in_reg7_5, in_reg7_6, in_reg7_7, in_reg8_0, in_reg8_1, in_reg8_2, in_reg8_3, in_reg8_4, in_reg8_5, in_reg8_6, in_reg8_7, in_reg8_8, in_reg9_0, in_reg9_1, in_reg9_2, in_reg9_3, in_reg9_4, in_reg9_5, in_reg9_6, in_reg9_7, in_reg9_8, in_reg9_9, in_reg10_0, in_reg10_1, in_reg10_2, in_reg10_3, in_reg10_4, in_reg10_5, in_reg10_6, in_reg10_7, in_reg10_8, in_reg10_9, in_reg10_10, in_reg11_0, in_reg11_1, in_reg11_2, in_reg11_3, in_reg11_4, in_reg11_5, in_reg11_6, in_reg11_7, in_reg11_8, in_reg11_9, in_reg11_10, in_reg11_11, in_reg12_0, in_reg12_1, in_reg12_2, in_reg12_3, in_reg12_4, in_reg12_5, in_reg12_6, in_reg12_7, in_reg12_8, in_reg12_9, in_reg12_10, in_reg12_11, in_reg12_12, in_reg13_0, in_reg13_1, in_reg13_2, in_reg13_3, in_reg13_4, in_reg13_5, in_reg13_6, in_reg13_7, in_reg13_8, in_reg13_9, in_reg13_10, in_reg13_11, in_reg13_12, in_reg13_13, in_reg14_0, in_reg14_1, in_reg14_2, in_reg14_3, in_reg14_4, in_reg14_5, in_reg14_6, in_reg14_7, in_reg14_8, in_reg14_9, in_reg14_10, in_reg14_11, in_reg14_12, in_reg14_13, in_reg14_14, in_reg15_0, in_reg15_1, in_reg15_2, in_reg15_3, in_reg15_4, in_reg15_5, in_reg15_6, in_reg15_7, in_reg15_8, in_reg15_9, in_reg15_10, in_reg15_11, in_reg15_12, in_reg15_13, in_reg15_14, in_reg15_15;

reg [31:0] in_pre_reg_0, in_pre_reg_1, in_pre_reg_2;

always @(posedge clk) begin
	if (command == 2'b01)
	begin
	case(col)
		2'd0: in_pre_reg_0 <= input0;
		2'd1: in_pre_reg_1 <= input0;
		2'd2: in_pre_reg_2 <= input0;
		default:;
	endcase
	end
	else
	begin
		in_pre_reg_0 <= in_pre_reg_0;
		in_pre_reg_1 <= in_pre_reg_1;
		in_pre_reg_2 <= in_pre_reg_2;
	end
	
end

assign fifo_enable = (col ==2'b11) && (command == 2'b10);

always@ (posedge clk)
begin
	if (fifo_enable)
	begin
		in_reg0_0 <= in_pre_reg_0[7:0];
		in_reg1_0 <= in_pre_reg_0[15:8];
		in_reg2_0 <= in_pre_reg_0[23:16];
		in_reg3_0 <= in_pre_reg_0[31:24];
		in_reg4_0 <= in_pre_reg_1[7:0];
		in_reg5_0 <= in_pre_reg_1[15:8];
		in_reg6_0 <= in_pre_reg_1[23:16];
		in_reg7_0 <= in_pre_reg_1[31:24];
		in_reg8_0 <= in_pre_reg_2[7:0];
		in_reg9_0 <= in_pre_reg_2[15:8];
		in_reg10_0 <= in_pre_reg_2[23:16];
		in_reg11_0 <= in_pre_reg_2[31:24];
		in_reg12_0 <= input0[7:0];
		in_reg13_0 <= input0[15:8];
		in_reg14_0 <= input0[23:16];
		in_reg15_0 <= input0[31:24];
		
		in_reg1_1 <= in_reg1_0;
		in_reg2_1 <= in_reg2_0;
		in_reg2_2 <= in_reg2_1;
		in_reg3_1 <= in_reg3_0;
		in_reg3_2 <= in_reg3_1;
		in_reg3_3 <= in_reg3_2;
		in_reg4_1 <= in_reg4_0;
		in_reg4_2 <= in_reg4_1;
		in_reg4_3 <= in_reg4_2;
		in_reg4_4 <= in_reg4_3;
		in_reg5_1 <= in_reg5_0;
		in_reg5_2 <= in_reg5_1;
		in_reg5_3 <= in_reg5_2;
		in_reg5_4 <= in_reg5_3;
		in_reg5_5 <= in_reg5_4;
		in_reg6_1 <= in_reg6_0;
		in_reg6_2 <= in_reg6_1;
		in_reg6_3 <= in_reg6_2;
		in_reg6_4 <= in_reg6_3;
		in_reg6_5 <= in_reg6_4;
		in_reg6_6 <= in_reg6_5;
		in_reg7_1 <= in_reg7_0;
		in_reg7_2 <= in_reg7_1;
		in_reg7_3 <= in_reg7_2;
		in_reg7_4 <= in_reg7_3;
		in_reg7_5 <= in_reg7_4;
		in_reg7_6 <= in_reg7_5;
		in_reg7_7 <= in_reg7_6;
		in_reg8_1 <= in_reg8_0;
		in_reg8_2 <= in_reg8_1;
		in_reg8_3 <= in_reg8_2;
		in_reg8_4 <= in_reg8_3;
		in_reg8_5 <= in_reg8_4;
		in_reg8_6 <= in_reg8_5;
		in_reg8_7 <= in_reg8_6;
		in_reg8_8 <= in_reg8_7;
		in_reg9_1 <= in_reg9_0;
		in_reg9_2 <= in_reg9_1;
		in_reg9_3 <= in_reg9_2;
		in_reg9_4 <= in_reg9_3;
		in_reg9_5 <= in_reg9_4;
		in_reg9_6 <= in_reg9_5;
		in_reg9_7 <= in_reg9_6;
		in_reg9_8 <= in_reg9_7;
		in_reg9_9 <= in_reg9_8;
		in_reg10_1 <= in_reg10_0;
		in_reg10_2 <= in_reg10_1;
		in_reg10_3 <= in_reg10_2;
		in_reg10_4 <= in_reg10_3;
		in_reg10_5 <= in_reg10_4;
		in_reg10_6 <= in_reg10_5;
		in_reg10_7 <= in_reg10_6;
		in_reg10_8 <= in_reg10_7;
		in_reg10_9 <= in_reg10_8;
		in_reg10_10 <= in_reg10_9;
		in_reg11_1 <= in_reg11_0;
		in_reg11_2 <= in_reg11_1;
		in_reg11_3 <= in_reg11_2;
		in_reg11_4 <= in_reg11_3;
		in_reg11_5 <= in_reg11_4;
		in_reg11_6 <= in_reg11_5;
		in_reg11_7 <= in_reg11_6;
		in_reg11_8 <= in_reg11_7;
		in_reg11_9 <= in_reg11_8;
		in_reg11_10 <= in_reg11_9;
		in_reg11_11 <= in_reg11_10;
		in_reg12_1 <= in_reg12_0;
		in_reg12_2 <= in_reg12_1;
		in_reg12_3 <= in_reg12_2;
		in_reg12_4 <= in_reg12_3;
		in_reg12_5 <= in_reg12_4;
		in_reg12_6 <= in_reg12_5;
		in_reg12_7 <= in_reg12_6;
		in_reg12_8 <= in_reg12_7;
		in_reg12_9 <= in_reg12_8;
		in_reg12_10 <= in_reg12_9;
		in_reg12_11 <= in_reg12_10;
		in_reg12_12 <= in_reg12_11;
		in_reg13_1 <= in_reg13_0;
		in_reg13_2 <= in_reg13_1;
		in_reg13_3 <= in_reg13_2;
		in_reg13_4 <= in_reg13_3;
		in_reg13_5 <= in_reg13_4;
		in_reg13_6 <= in_reg13_5;
		in_reg13_7 <= in_reg13_6;
		in_reg13_8 <= in_reg13_7;
		in_reg13_9 <= in_reg13_8;
		in_reg13_10 <= in_reg13_9;
		in_reg13_11 <= in_reg13_10;
		in_reg13_12 <= in_reg13_11;
		in_reg13_13 <= in_reg13_12;
		in_reg14_1 <= in_reg14_0;
		in_reg14_2 <= in_reg14_1;
		in_reg14_3 <= in_reg14_2;
		in_reg14_4 <= in_reg14_3;
		in_reg14_5 <= in_reg14_4;
		in_reg14_6 <= in_reg14_5;
		in_reg14_7 <= in_reg14_6;
		in_reg14_8 <= in_reg14_7;
		in_reg14_9 <= in_reg14_8;
		in_reg14_10 <= in_reg14_9;
		in_reg14_11 <= in_reg14_10;
		in_reg14_12 <= in_reg14_11;
		in_reg14_13 <= in_reg14_12;
		in_reg14_14 <= in_reg14_13;
		in_reg15_1 <= in_reg15_0;
		in_reg15_2 <= in_reg15_1;
		in_reg15_3 <= in_reg15_2;
		in_reg15_4 <= in_reg15_3;
		in_reg15_5 <= in_reg15_4;
		in_reg15_6 <= in_reg15_5;
		in_reg15_7 <= in_reg15_6;
		in_reg15_8 <= in_reg15_7;
		in_reg15_9 <= in_reg15_8;
		in_reg15_10 <= in_reg15_9;
		in_reg15_11 <= in_reg15_10;
		in_reg15_12 <= in_reg15_11;
		in_reg15_13 <= in_reg15_12;
		in_reg15_14 <= in_reg15_13;
		in_reg15_15 <= in_reg15_14;
		
	end
	else
	begin
		in_reg0_0 <= in_reg0_0;
		in_reg1_0 <= in_reg1_0;
		in_reg1_1 <= in_reg1_1;
		in_reg2_0 <= in_reg2_0;
		in_reg2_1 <= in_reg2_1;
		in_reg2_2 <= in_reg2_2;
		in_reg3_0 <= in_reg3_0;
		in_reg3_1 <= in_reg3_1;
		in_reg3_2 <= in_reg3_2;
		in_reg3_3 <= in_reg3_3;
		in_reg4_0 <= in_reg4_0;
		in_reg4_1 <= in_reg4_1;
		in_reg4_2 <= in_reg4_2;
		in_reg4_3 <= in_reg4_3;
		in_reg4_4 <= in_reg4_4;
		in_reg5_0 <= in_reg5_0;
		in_reg5_1 <= in_reg5_1;
		in_reg5_2 <= in_reg5_2;
		in_reg5_3 <= in_reg5_3;
		in_reg5_4 <= in_reg5_4;
		in_reg5_5 <= in_reg5_5;
		in_reg6_0 <= in_reg6_0;
		in_reg6_1 <= in_reg6_1;
		in_reg6_2 <= in_reg6_2;
		in_reg6_3 <= in_reg6_3;
		in_reg6_4 <= in_reg6_4;
		in_reg6_5 <= in_reg6_5;
		in_reg6_6 <= in_reg6_6;
		in_reg7_0 <= in_reg7_0;
		in_reg7_1 <= in_reg7_1;
		in_reg7_2 <= in_reg7_2;
		in_reg7_3 <= in_reg7_3;
		in_reg7_4 <= in_reg7_4;
		in_reg7_5 <= in_reg7_5;
		in_reg7_6 <= in_reg7_6;
		in_reg7_7 <= in_reg7_7;
		in_reg8_0 <= in_reg8_0;
		in_reg8_1 <= in_reg8_1;
		in_reg8_2 <= in_reg8_2;
		in_reg8_3 <= in_reg8_3;
		in_reg8_4 <= in_reg8_4;
		in_reg8_5 <= in_reg8_5;
		in_reg8_6 <= in_reg8_6;
		in_reg8_7 <= in_reg8_7;
		in_reg8_8 <= in_reg8_8;
		in_reg9_0 <= in_reg9_0;
		in_reg9_1 <= in_reg9_1;
		in_reg9_2 <= in_reg9_2;
		in_reg9_3 <= in_reg9_3;
		in_reg9_4 <= in_reg9_4;
		in_reg9_5 <= in_reg9_5;
		in_reg9_6 <= in_reg9_6;
		in_reg9_7 <= in_reg9_7;
		in_reg9_8 <= in_reg9_8;
		in_reg9_9 <= in_reg9_9;
		in_reg10_0 <= in_reg10_0;
		in_reg10_1 <= in_reg10_1;
		in_reg10_2 <= in_reg10_2;
		in_reg10_3 <= in_reg10_3;
		in_reg10_4 <= in_reg10_4;
		in_reg10_5 <= in_reg10_5;
		in_reg10_6 <= in_reg10_6;
		in_reg10_7 <= in_reg10_7;
		in_reg10_8 <= in_reg10_8;
		in_reg10_9 <= in_reg10_9;
		in_reg10_10 <= in_reg10_10;
		in_reg11_0 <= in_reg11_0;
		in_reg11_1 <= in_reg11_1;
		in_reg11_2 <= in_reg11_2;
		in_reg11_3 <= in_reg11_3;
		in_reg11_4 <= in_reg11_4;
		in_reg11_5 <= in_reg11_5;
		in_reg11_6 <= in_reg11_6;
		in_reg11_7 <= in_reg11_7;
		in_reg11_8 <= in_reg11_8;
		in_reg11_9 <= in_reg11_9;
		in_reg11_10 <= in_reg11_10;
		in_reg11_11 <= in_reg11_11;
		in_reg12_0 <= in_reg12_0;
		in_reg12_1 <= in_reg12_1;
		in_reg12_2 <= in_reg12_2;
		in_reg12_3 <= in_reg12_3;
		in_reg12_4 <= in_reg12_4;
		in_reg12_5 <= in_reg12_5;
		in_reg12_6 <= in_reg12_6;
		in_reg12_7 <= in_reg12_7;
		in_reg12_8 <= in_reg12_8;
		in_reg12_9 <= in_reg12_9;
		in_reg12_10 <= in_reg12_10;
		in_reg12_11 <= in_reg12_11;
		in_reg12_12 <= in_reg12_12;
		in_reg13_0 <= in_reg13_0;
		in_reg13_1 <= in_reg13_1;
		in_reg13_2 <= in_reg13_2;
		in_reg13_3 <= in_reg13_3;
		in_reg13_4 <= in_reg13_4;
		in_reg13_5 <= in_reg13_5;
		in_reg13_6 <= in_reg13_6;
		in_reg13_7 <= in_reg13_7;
		in_reg13_8 <= in_reg13_8;
		in_reg13_9 <= in_reg13_9;
		in_reg13_10 <= in_reg13_10;
		in_reg13_11 <= in_reg13_11;
		in_reg13_12 <= in_reg13_12;
		in_reg13_13 <= in_reg13_13;
		in_reg14_0 <= in_reg14_0;
		in_reg14_1 <= in_reg14_1;
		in_reg14_2 <= in_reg14_2;
		in_reg14_3 <= in_reg14_3;
		in_reg14_4 <= in_reg14_4;
		in_reg14_5 <= in_reg14_5;
		in_reg14_6 <= in_reg14_6;
		in_reg14_7 <= in_reg14_7;
		in_reg14_8 <= in_reg14_8;
		in_reg14_9 <= in_reg14_9;
		in_reg14_10 <= in_reg14_10;
		in_reg14_11 <= in_reg14_11;
		in_reg14_12 <= in_reg14_12;
		in_reg14_13 <= in_reg14_13;
		in_reg14_14 <= in_reg14_14;
		in_reg15_0 <= in_reg15_0;
		in_reg15_1 <= in_reg15_1;
		in_reg15_2 <= in_reg15_2;
		in_reg15_3 <= in_reg15_3;
		in_reg15_4 <= in_reg15_4;
		in_reg15_5 <= in_reg15_5;
		in_reg15_6 <= in_reg15_6;
		in_reg15_7 <= in_reg15_7;
		in_reg15_8 <= in_reg15_8;
		in_reg15_9 <= in_reg15_9;
		in_reg15_10 <= in_reg15_10;
		in_reg15_11 <= in_reg15_11;
		in_reg15_12 <= in_reg15_12;
		in_reg15_13 <= in_reg15_13;
		in_reg15_14 <= in_reg15_14;
		in_reg15_15 <= in_reg15_15;	
	end
end

assign output0 = in_reg0_0;
assign output1 = in_reg1_1;
assign output2 = in_reg2_2;
assign output3 = in_reg3_3;
assign output4 = in_reg4_4;
assign output5 = in_reg5_5;
assign output6 = in_reg6_6;
assign output7 = in_reg7_7;
assign output8 = in_reg8_8;
assign output9 = in_reg9_9;
assign output10 = in_reg10_10;
assign output11 = in_reg11_11;
assign output12 = in_reg12_12;
assign output13 = in_reg13_13;
assign output14 = in_reg14_14;
assign output15 = in_reg15_15;


endmodule 
