module SA(w_input, input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15,
output0, output1, output2, output3, output4, output5, output6, output7, output8, output9, output10, output11, output12, output13, output14, output15, 
command, col, resetn,clk);
input [31:0] w_input;
input signed [7:0] input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15;
input [1:0] command;
input [1:0] col;
output signed [7:0] output0, output1, output2, output3, output4, output5, output6, output7, output8, output9, output10, output11, output12, output13, output14, output15;
input clk , resetn;

wire load_enable;
reg [31:0]  weight_reg00, weight_reg01, weight_reg02, weight_reg03, weight_reg10, weight_reg11, weight_reg12, weight_reg13, weight_reg20, weight_reg21, weight_reg22, weight_reg23, weight_reg30, weight_reg31, weight_reg32, weight_reg33, weight_reg40, weight_reg41, weight_reg42, weight_reg43, weight_reg50, weight_reg51, weight_reg52, weight_reg53, weight_reg60, weight_reg61, weight_reg62, weight_reg63, weight_reg70, weight_reg71, weight_reg72, weight_reg73, weight_reg80, weight_reg81, weight_reg82, weight_reg83, weight_reg90, weight_reg91, weight_reg92, weight_reg93, weight_reg100, weight_reg101, weight_reg102, weight_reg103, weight_reg110, weight_reg111, weight_reg112, weight_reg113, weight_reg120, weight_reg121, weight_reg122, weight_reg123, weight_reg130, weight_reg131, weight_reg132, weight_reg133, weight_reg140, weight_reg141, weight_reg142, weight_reg143, weight_reg150, weight_reg151, weight_reg152, weight_reg153;

reg [31:0] weight_pre_reg_0, weight_pre_reg_1, weight_pre_reg_2;

always @(posedge clk) begin
	if (command == 2'b00)
	begin
	case(col)
		2'd0: weight_pre_reg_0 <= w_input;
		2'd1: weight_pre_reg_1 <= w_input;
		2'd2: weight_pre_reg_2 <= w_input;
		default:;
	endcase
	end
	else
	begin
		weight_pre_reg_0 <= weight_pre_reg_0;
		weight_pre_reg_1 <= weight_pre_reg_1;
		weight_pre_reg_2 <= weight_pre_reg_2;
	end
	
end

assign load_enable = (col ==2'b11) && (command == 2'b00);

always@ (posedge clk)
begin
	if (load_enable)
	begin
		weight_reg00 <= weight_pre_reg_0;
		weight_reg01 <= weight_pre_reg_1;
		weight_reg02 <= weight_pre_reg_2;
		weight_reg03 <= w_input;
		
		weight_reg10 <= weight_reg00;
		weight_reg20 <= weight_reg10;
		weight_reg30 <= weight_reg20;
		weight_reg40 <= weight_reg30;
		weight_reg50 <= weight_reg40;
		weight_reg60 <= weight_reg50;
		weight_reg70 <= weight_reg60;
		weight_reg80 <= weight_reg70;
		weight_reg90 <= weight_reg80;
		weight_reg100 <= weight_reg90;
		weight_reg110 <= weight_reg100;
		weight_reg120 <= weight_reg110;
		weight_reg130 <= weight_reg120;
		weight_reg140 <= weight_reg130;
		weight_reg150 <= weight_reg140;
		weight_reg11 <= weight_reg01;
		weight_reg21 <= weight_reg11;
		weight_reg31 <= weight_reg21;
		weight_reg41 <= weight_reg31;
		weight_reg51 <= weight_reg41;
		weight_reg61 <= weight_reg51;
		weight_reg71 <= weight_reg61;
		weight_reg81 <= weight_reg71;
		weight_reg91 <= weight_reg81;
		weight_reg101 <= weight_reg91;
		weight_reg111 <= weight_reg101;
		weight_reg121 <= weight_reg111;
		weight_reg131 <= weight_reg121;
		weight_reg141 <= weight_reg131;
		weight_reg151 <= weight_reg141;
		weight_reg12 <= weight_reg02;
		weight_reg22 <= weight_reg12;
		weight_reg32 <= weight_reg22;
		weight_reg42 <= weight_reg32;
		weight_reg52 <= weight_reg42;
		weight_reg62 <= weight_reg52;
		weight_reg72 <= weight_reg62;
		weight_reg82 <= weight_reg72;
		weight_reg92 <= weight_reg82;
		weight_reg102 <= weight_reg92;
		weight_reg112 <= weight_reg102;
		weight_reg122 <= weight_reg112;
		weight_reg132 <= weight_reg122;
		weight_reg142 <= weight_reg132;
		weight_reg152 <= weight_reg142;
		weight_reg13 <= weight_reg03;
		weight_reg23 <= weight_reg13;
		weight_reg33 <= weight_reg23;
		weight_reg43 <= weight_reg33;
		weight_reg53 <= weight_reg43;
		weight_reg63 <= weight_reg53;
		weight_reg73 <= weight_reg63;
		weight_reg83 <= weight_reg73;
		weight_reg93 <= weight_reg83;
		weight_reg103 <= weight_reg93;
		weight_reg113 <= weight_reg103;
		weight_reg123 <= weight_reg113;
		weight_reg133 <= weight_reg123;
		weight_reg143 <= weight_reg133;
		weight_reg153 <= weight_reg143;
	end
end

reg signed [7:0] in_reg0_0, in_reg0_1, in_reg0_2, in_reg0_3, in_reg0_4, in_reg0_5, in_reg0_6, in_reg0_7, in_reg0_8, in_reg0_9, in_reg0_10, in_reg0_11, in_reg0_12, in_reg0_13, in_reg0_14, in_reg0_15, in_reg1_0, in_reg1_1, in_reg1_2, in_reg1_3, in_reg1_4, in_reg1_5, in_reg1_6, in_reg1_7, in_reg1_8, in_reg1_9, in_reg1_10, in_reg1_11, in_reg1_12, in_reg1_13, in_reg1_14, in_reg1_15, in_reg2_0, in_reg2_1, in_reg2_2, in_reg2_3, in_reg2_4, in_reg2_5, in_reg2_6, in_reg2_7, in_reg2_8, in_reg2_9, in_reg2_10, in_reg2_11, in_reg2_12, in_reg2_13, in_reg2_14, in_reg2_15, in_reg3_0, in_reg3_1, in_reg3_2, in_reg3_3, in_reg3_4, in_reg3_5, in_reg3_6, in_reg3_7, in_reg3_8, in_reg3_9, in_reg3_10, in_reg3_11, in_reg3_12, in_reg3_13, in_reg3_14, in_reg3_15, in_reg4_0, in_reg4_1, in_reg4_2, in_reg4_3, in_reg4_4, in_reg4_5, in_reg4_6, in_reg4_7, in_reg4_8, in_reg4_9, in_reg4_10, in_reg4_11, in_reg4_12, in_reg4_13, in_reg4_14, in_reg4_15, in_reg5_0, in_reg5_1, in_reg5_2, in_reg5_3, in_reg5_4, in_reg5_5, in_reg5_6, in_reg5_7, in_reg5_8, in_reg5_9, in_reg5_10, in_reg5_11, in_reg5_12, in_reg5_13, in_reg5_14, in_reg5_15, in_reg6_0, in_reg6_1, in_reg6_2, in_reg6_3, in_reg6_4, in_reg6_5, in_reg6_6, in_reg6_7, in_reg6_8, in_reg6_9, in_reg6_10, in_reg6_11, in_reg6_12, in_reg6_13, in_reg6_14, in_reg6_15, in_reg7_0, in_reg7_1, in_reg7_2, in_reg7_3, in_reg7_4, in_reg7_5, in_reg7_6, in_reg7_7, in_reg7_8, in_reg7_9, in_reg7_10, in_reg7_11, in_reg7_12, in_reg7_13, in_reg7_14, in_reg7_15, in_reg8_0, in_reg8_1, in_reg8_2, in_reg8_3, in_reg8_4, in_reg8_5, in_reg8_6, in_reg8_7, in_reg8_8, in_reg8_9, in_reg8_10, in_reg8_11, in_reg8_12, in_reg8_13, in_reg8_14, in_reg8_15, in_reg9_0, in_reg9_1, in_reg9_2, in_reg9_3, in_reg9_4, in_reg9_5, in_reg9_6, in_reg9_7, in_reg9_8, in_reg9_9, in_reg9_10, in_reg9_11, in_reg9_12, in_reg9_13, in_reg9_14, in_reg9_15, in_reg10_0, in_reg10_1, in_reg10_2, in_reg10_3, in_reg10_4, in_reg10_5, in_reg10_6, in_reg10_7, in_reg10_8, in_reg10_9, in_reg10_10, in_reg10_11, in_reg10_12, in_reg10_13, in_reg10_14, in_reg10_15, in_reg11_0, in_reg11_1, in_reg11_2, in_reg11_3, in_reg11_4, in_reg11_5, in_reg11_6, in_reg11_7, in_reg11_8, in_reg11_9, in_reg11_10, in_reg11_11, in_reg11_12, in_reg11_13, in_reg11_14, in_reg11_15, in_reg12_0, in_reg12_1, in_reg12_2, in_reg12_3, in_reg12_4, in_reg12_5, in_reg12_6, in_reg12_7, in_reg12_8, in_reg12_9, in_reg12_10, in_reg12_11, in_reg12_12, in_reg12_13, in_reg12_14, in_reg12_15, in_reg13_0, in_reg13_1, in_reg13_2, in_reg13_3, in_reg13_4, in_reg13_5, in_reg13_6, in_reg13_7, in_reg13_8, in_reg13_9, in_reg13_10, in_reg13_11, in_reg13_12, in_reg13_13, in_reg13_14, in_reg13_15, in_reg14_0, in_reg14_1, in_reg14_2, in_reg14_3, in_reg14_4, in_reg14_5, in_reg14_6, in_reg14_7, in_reg14_8, in_reg14_9, in_reg14_10, in_reg14_11, in_reg14_12, in_reg14_13, in_reg14_14, in_reg14_15, in_reg15_0, in_reg15_1, in_reg15_2, in_reg15_3, in_reg15_4, in_reg15_5, in_reg15_6, in_reg15_7, in_reg15_8, in_reg15_9, in_reg15_10, in_reg15_11, in_reg15_12, in_reg15_13, in_reg15_14, in_reg15_15;

reg signed [7:0] acc_reg0_0, acc_reg0_1, acc_reg0_2, acc_reg0_3, acc_reg0_4, acc_reg0_5, acc_reg0_6, acc_reg0_7, acc_reg0_8, acc_reg0_9, acc_reg0_10, acc_reg0_11, acc_reg0_12, acc_reg0_13, acc_reg0_14, acc_reg0_15, acc_reg1_0, acc_reg1_1, acc_reg1_2, acc_reg1_3, acc_reg1_4, acc_reg1_5, acc_reg1_6, acc_reg1_7, acc_reg1_8, acc_reg1_9, acc_reg1_10, acc_reg1_11, acc_reg1_12, acc_reg1_13, acc_reg1_14, acc_reg1_15, acc_reg2_0, acc_reg2_1, acc_reg2_2, acc_reg2_3, acc_reg2_4, acc_reg2_5, acc_reg2_6, acc_reg2_7, acc_reg2_8, acc_reg2_9, acc_reg2_10, acc_reg2_11, acc_reg2_12, acc_reg2_13, acc_reg2_14, acc_reg2_15, acc_reg3_0, acc_reg3_1, acc_reg3_2, acc_reg3_3, acc_reg3_4, acc_reg3_5, acc_reg3_6, acc_reg3_7, acc_reg3_8, acc_reg3_9, acc_reg3_10, acc_reg3_11, acc_reg3_12, acc_reg3_13, acc_reg3_14, acc_reg3_15, acc_reg4_0, acc_reg4_1, acc_reg4_2, acc_reg4_3, acc_reg4_4, acc_reg4_5, acc_reg4_6, acc_reg4_7, acc_reg4_8, acc_reg4_9, acc_reg4_10, acc_reg4_11, acc_reg4_12, acc_reg4_13, acc_reg4_14, acc_reg4_15, acc_reg5_0, acc_reg5_1, acc_reg5_2, acc_reg5_3, acc_reg5_4, acc_reg5_5, acc_reg5_6, acc_reg5_7, acc_reg5_8, acc_reg5_9, acc_reg5_10, acc_reg5_11, acc_reg5_12, acc_reg5_13, acc_reg5_14, acc_reg5_15, acc_reg6_0, acc_reg6_1, acc_reg6_2, acc_reg6_3, acc_reg6_4, acc_reg6_5, acc_reg6_6, acc_reg6_7, acc_reg6_8, acc_reg6_9, acc_reg6_10, acc_reg6_11, acc_reg6_12, acc_reg6_13, acc_reg6_14, acc_reg6_15, acc_reg7_0, acc_reg7_1, acc_reg7_2, acc_reg7_3, acc_reg7_4, acc_reg7_5, acc_reg7_6, acc_reg7_7, acc_reg7_8, acc_reg7_9, acc_reg7_10, acc_reg7_11, acc_reg7_12, acc_reg7_13, acc_reg7_14, acc_reg7_15, acc_reg8_0, acc_reg8_1, acc_reg8_2, acc_reg8_3, acc_reg8_4, acc_reg8_5, acc_reg8_6, acc_reg8_7, acc_reg8_8, acc_reg8_9, acc_reg8_10, acc_reg8_11, acc_reg8_12, acc_reg8_13, acc_reg8_14, acc_reg8_15, acc_reg9_0, acc_reg9_1, acc_reg9_2, acc_reg9_3, acc_reg9_4, acc_reg9_5, acc_reg9_6, acc_reg9_7, acc_reg9_8, acc_reg9_9, acc_reg9_10, acc_reg9_11, acc_reg9_12, acc_reg9_13, acc_reg9_14, acc_reg9_15, acc_reg10_0, acc_reg10_1, acc_reg10_2, acc_reg10_3, acc_reg10_4, acc_reg10_5, acc_reg10_6, acc_reg10_7, acc_reg10_8, acc_reg10_9, acc_reg10_10, acc_reg10_11, acc_reg10_12, acc_reg10_13, acc_reg10_14, acc_reg10_15, acc_reg11_0, acc_reg11_1, acc_reg11_2, acc_reg11_3, acc_reg11_4, acc_reg11_5, acc_reg11_6, acc_reg11_7, acc_reg11_8, acc_reg11_9, acc_reg11_10, acc_reg11_11, acc_reg11_12, acc_reg11_13, acc_reg11_14, acc_reg11_15, acc_reg12_0, acc_reg12_1, acc_reg12_2, acc_reg12_3, acc_reg12_4, acc_reg12_5, acc_reg12_6, acc_reg12_7, acc_reg12_8, acc_reg12_9, acc_reg12_10, acc_reg12_11, acc_reg12_12, acc_reg12_13, acc_reg12_14, acc_reg12_15, acc_reg13_0, acc_reg13_1, acc_reg13_2, acc_reg13_3, acc_reg13_4, acc_reg13_5, acc_reg13_6, acc_reg13_7, acc_reg13_8, acc_reg13_9, acc_reg13_10, acc_reg13_11, acc_reg13_12, acc_reg13_13, acc_reg13_14, acc_reg13_15, acc_reg14_0, acc_reg14_1, acc_reg14_2, acc_reg14_3, acc_reg14_4, acc_reg14_5, acc_reg14_6, acc_reg14_7, acc_reg14_8, acc_reg14_9, acc_reg14_10, acc_reg14_11, acc_reg14_12, acc_reg14_13, acc_reg14_14, acc_reg14_15, acc_reg15_0, acc_reg15_1, acc_reg15_2, acc_reg15_3, acc_reg15_4, acc_reg15_5, acc_reg15_6, acc_reg15_7, acc_reg15_8, acc_reg15_9, acc_reg15_10, acc_reg15_11, acc_reg15_12, acc_reg15_13, acc_reg15_14, acc_reg15_15;


wire signed [7:0] acc_wire0_0, acc_wire0_1, acc_wire0_2, acc_wire0_3, acc_wire0_4, acc_wire0_5, acc_wire0_6, acc_wire0_7, acc_wire0_8, acc_wire0_9, acc_wire0_10, acc_wire0_11, acc_wire0_12, acc_wire0_13, acc_wire0_14, acc_wire0_15, acc_wire1_0, acc_wire1_1, acc_wire1_2, acc_wire1_3, acc_wire1_4, acc_wire1_5, acc_wire1_6, acc_wire1_7, acc_wire1_8, acc_wire1_9, acc_wire1_10, acc_wire1_11, acc_wire1_12, acc_wire1_13, acc_wire1_14, acc_wire1_15, acc_wire2_0, acc_wire2_1, acc_wire2_2, acc_wire2_3, acc_wire2_4, acc_wire2_5, acc_wire2_6, acc_wire2_7, acc_wire2_8, acc_wire2_9, acc_wire2_10, acc_wire2_11, acc_wire2_12, acc_wire2_13, acc_wire2_14, acc_wire2_15, acc_wire3_0, acc_wire3_1, acc_wire3_2, acc_wire3_3, acc_wire3_4, acc_wire3_5, acc_wire3_6, acc_wire3_7, acc_wire3_8, acc_wire3_9, acc_wire3_10, acc_wire3_11, acc_wire3_12, acc_wire3_13, acc_wire3_14, acc_wire3_15, acc_wire4_0, acc_wire4_1, acc_wire4_2, acc_wire4_3, acc_wire4_4, acc_wire4_5, acc_wire4_6, acc_wire4_7, acc_wire4_8, acc_wire4_9, acc_wire4_10, acc_wire4_11, acc_wire4_12, acc_wire4_13, acc_wire4_14, acc_wire4_15, acc_wire5_0, acc_wire5_1, acc_wire5_2, acc_wire5_3, acc_wire5_4, acc_wire5_5, acc_wire5_6, acc_wire5_7, acc_wire5_8, acc_wire5_9, acc_wire5_10, acc_wire5_11, acc_wire5_12, acc_wire5_13, acc_wire5_14, acc_wire5_15, acc_wire6_0, acc_wire6_1, acc_wire6_2, acc_wire6_3, acc_wire6_4, acc_wire6_5, acc_wire6_6, acc_wire6_7, acc_wire6_8, acc_wire6_9, acc_wire6_10, acc_wire6_11, acc_wire6_12, acc_wire6_13, acc_wire6_14, acc_wire6_15, acc_wire7_0, acc_wire7_1, acc_wire7_2, acc_wire7_3, acc_wire7_4, acc_wire7_5, acc_wire7_6, acc_wire7_7, acc_wire7_8, acc_wire7_9, acc_wire7_10, acc_wire7_11, acc_wire7_12, acc_wire7_13, acc_wire7_14, acc_wire7_15, acc_wire8_0, acc_wire8_1, acc_wire8_2, acc_wire8_3, acc_wire8_4, acc_wire8_5, acc_wire8_6, acc_wire8_7, acc_wire8_8, acc_wire8_9, acc_wire8_10, acc_wire8_11, acc_wire8_12, acc_wire8_13, acc_wire8_14, acc_wire8_15, acc_wire9_0, acc_wire9_1, acc_wire9_2, acc_wire9_3, acc_wire9_4, acc_wire9_5, acc_wire9_6, acc_wire9_7, acc_wire9_8, acc_wire9_9, acc_wire9_10, acc_wire9_11, acc_wire9_12, acc_wire9_13, acc_wire9_14, acc_wire9_15, acc_wire10_0, acc_wire10_1, acc_wire10_2, acc_wire10_3, acc_wire10_4, acc_wire10_5, acc_wire10_6, acc_wire10_7, acc_wire10_8, acc_wire10_9, acc_wire10_10, acc_wire10_11, acc_wire10_12, acc_wire10_13, acc_wire10_14, acc_wire10_15, acc_wire11_0, acc_wire11_1, acc_wire11_2, acc_wire11_3, acc_wire11_4, acc_wire11_5, acc_wire11_6, acc_wire11_7, acc_wire11_8, acc_wire11_9, acc_wire11_10, acc_wire11_11, acc_wire11_12, acc_wire11_13, acc_wire11_14, acc_wire11_15, acc_wire12_0, acc_wire12_1, acc_wire12_2, acc_wire12_3, acc_wire12_4, acc_wire12_5, acc_wire12_6, acc_wire12_7, acc_wire12_8, acc_wire12_9, acc_wire12_10, acc_wire12_11, acc_wire12_12, acc_wire12_13, acc_wire12_14, acc_wire12_15, acc_wire13_0, acc_wire13_1, acc_wire13_2, acc_wire13_3, acc_wire13_4, acc_wire13_5, acc_wire13_6, acc_wire13_7, acc_wire13_8, acc_wire13_9, acc_wire13_10, acc_wire13_11, acc_wire13_12, acc_wire13_13, acc_wire13_14, acc_wire13_15, acc_wire14_0, acc_wire14_1, acc_wire14_2, acc_wire14_3, acc_wire14_4, acc_wire14_5, acc_wire14_6, acc_wire14_7, acc_wire14_8, acc_wire14_9, acc_wire14_10, acc_wire14_11, acc_wire14_12, acc_wire14_13, acc_wire14_14, acc_wire14_15, acc_wire15_0, acc_wire15_1, acc_wire15_2, acc_wire15_3, acc_wire15_4, acc_wire15_5, acc_wire15_6, acc_wire15_7, acc_wire15_8, acc_wire15_9, acc_wire15_10, acc_wire15_11, acc_wire15_12, acc_wire15_13, acc_wire15_14, acc_wire15_15;

PE PE0_0(.in(input0), .acc(8'b0), .w(weight_reg00[7:0]), .out(acc_wire0_0), .resetn(resetn),.clk(clk));
PE PE0_1(.in(in_reg0_1), .acc(8'b0), .w(weight_reg00[15:8]), .out(acc_wire0_1), .resetn(resetn),.clk(clk));
PE PE0_2(.in(in_reg0_2), .acc(8'b0), .w(weight_reg00[23:16]), .out(acc_wire0_2), .resetn(resetn),.clk(clk));
PE PE0_3(.in(in_reg0_3), .acc(8'b0), .w(weight_reg00[31:24]), .out(acc_wire0_3), .resetn(resetn),.clk(clk));
PE PE0_4(.in(in_reg0_4), .acc(8'b0), .w(weight_reg01[7:0]), .out(acc_wire0_4), .resetn(resetn),.clk(clk));
PE PE0_5(.in(in_reg0_5), .acc(8'b0), .w(weight_reg01[15:8]), .out(acc_wire0_5), .resetn(resetn),.clk(clk));
PE PE0_6(.in(in_reg0_6), .acc(8'b0), .w(weight_reg01[23:16]), .out(acc_wire0_6), .resetn(resetn),.clk(clk));
PE PE0_7(.in(in_reg0_7), .acc(8'b0), .w(weight_reg01[31:24]), .out(acc_wire0_7), .resetn(resetn),.clk(clk));
PE PE0_8(.in(in_reg0_8), .acc(8'b0), .w(weight_reg02[7:0]), .out(acc_wire0_8), .resetn(resetn),.clk(clk));
PE PE0_9(.in(in_reg0_9), .acc(8'b0), .w(weight_reg02[15:8]), .out(acc_wire0_9), .resetn(resetn),.clk(clk));
PE PE0_10(.in(in_reg0_10), .acc(8'b0), .w(weight_reg02[23:16]), .out(acc_wire0_10), .resetn(resetn),.clk(clk));
PE PE0_11(.in(in_reg0_11), .acc(8'b0), .w(weight_reg02[31:24]), .out(acc_wire0_11), .resetn(resetn),.clk(clk));
PE PE0_12(.in(in_reg0_12), .acc(8'b0), .w(weight_reg03[7:0]), .out(acc_wire0_12), .resetn(resetn),.clk(clk));
PE PE0_13(.in(in_reg0_13), .acc(8'b0), .w(weight_reg03[15:8]), .out(acc_wire0_13), .resetn(resetn),.clk(clk));
PE PE0_14(.in(in_reg0_14), .acc(8'b0), .w(weight_reg03[23:16]), .out(acc_wire0_14), .resetn(resetn),.clk(clk));
PE PE0_15(.in(in_reg0_15), .acc(8'b0), .w(weight_reg03[31:24]), .out(acc_wire0_15), .resetn(resetn),.clk(clk));

PE PE1_0(.in(input1), .acc(acc_reg0_0), .w(weight_reg10[7:0]), .out(acc_wire1_0), .resetn(resetn),.clk(clk));
PE PE1_1(.in(in_reg1_1), .acc(acc_reg0_1), .w(weight_reg10[15:8]), .out(acc_wire1_1), .resetn(resetn),.clk(clk));
PE PE1_2(.in(in_reg1_2), .acc(acc_reg0_2), .w(weight_reg10[23:16]), .out(acc_wire1_2), .resetn(resetn),.clk(clk));
PE PE1_3(.in(in_reg1_3), .acc(acc_reg0_3), .w(weight_reg10[31:24]), .out(acc_wire1_3), .resetn(resetn),.clk(clk));
PE PE1_4(.in(in_reg1_4), .acc(acc_reg0_4), .w(weight_reg11[7:0]), .out(acc_wire1_4), .resetn(resetn),.clk(clk));
PE PE1_5(.in(in_reg1_5), .acc(acc_reg0_5), .w(weight_reg11[15:8]), .out(acc_wire1_5), .resetn(resetn),.clk(clk));
PE PE1_6(.in(in_reg1_6), .acc(acc_reg0_6), .w(weight_reg11[23:16]), .out(acc_wire1_6), .resetn(resetn),.clk(clk));
PE PE1_7(.in(in_reg1_7), .acc(acc_reg0_7), .w(weight_reg11[31:24]), .out(acc_wire1_7), .resetn(resetn),.clk(clk));
PE PE1_8(.in(in_reg1_8), .acc(acc_reg0_8), .w(weight_reg12[7:0]), .out(acc_wire1_8), .resetn(resetn),.clk(clk));
PE PE1_9(.in(in_reg1_9), .acc(acc_reg0_9), .w(weight_reg12[15:8]), .out(acc_wire1_9), .resetn(resetn),.clk(clk));
PE PE1_10(.in(in_reg1_10), .acc(acc_reg0_10), .w(weight_reg12[23:16]), .out(acc_wire1_10), .resetn(resetn),.clk(clk));
PE PE1_11(.in(in_reg1_11), .acc(acc_reg0_11), .w(weight_reg12[31:24]), .out(acc_wire1_11), .resetn(resetn),.clk(clk));
PE PE1_12(.in(in_reg1_12), .acc(acc_reg0_12), .w(weight_reg13[7:0]), .out(acc_wire1_12), .resetn(resetn),.clk(clk));
PE PE1_13(.in(in_reg1_13), .acc(acc_reg0_13), .w(weight_reg13[15:8]), .out(acc_wire1_13), .resetn(resetn),.clk(clk));
PE PE1_14(.in(in_reg1_14), .acc(acc_reg0_14), .w(weight_reg13[23:16]), .out(acc_wire1_14), .resetn(resetn),.clk(clk));
PE PE1_15(.in(in_reg1_15), .acc(acc_reg0_15), .w(weight_reg13[31:24]), .out(acc_wire1_15), .resetn(resetn),.clk(clk));

PE PE2_0(.in(input2), .acc(acc_reg1_0), .w(weight_reg20[7:0]), .out(acc_wire2_0), .resetn(resetn),.clk(clk));
PE PE2_1(.in(in_reg2_1), .acc(acc_reg1_1), .w(weight_reg20[15:8]), .out(acc_wire2_1), .resetn(resetn),.clk(clk));
PE PE2_2(.in(in_reg2_2), .acc(acc_reg1_2), .w(weight_reg20[23:16]), .out(acc_wire2_2), .resetn(resetn),.clk(clk));
PE PE2_3(.in(in_reg2_3), .acc(acc_reg1_3), .w(weight_reg20[31:24]), .out(acc_wire2_3), .resetn(resetn),.clk(clk));
PE PE2_4(.in(in_reg2_4), .acc(acc_reg1_4), .w(weight_reg21[7:0]), .out(acc_wire2_4), .resetn(resetn),.clk(clk));
PE PE2_5(.in(in_reg2_5), .acc(acc_reg1_5), .w(weight_reg21[15:8]), .out(acc_wire2_5), .resetn(resetn),.clk(clk));
PE PE2_6(.in(in_reg2_6), .acc(acc_reg1_6), .w(weight_reg21[23:16]), .out(acc_wire2_6), .resetn(resetn),.clk(clk));
PE PE2_7(.in(in_reg2_7), .acc(acc_reg1_7), .w(weight_reg21[31:24]), .out(acc_wire2_7), .resetn(resetn),.clk(clk));
PE PE2_8(.in(in_reg2_8), .acc(acc_reg1_8), .w(weight_reg22[7:0]), .out(acc_wire2_8), .resetn(resetn),.clk(clk));
PE PE2_9(.in(in_reg2_9), .acc(acc_reg1_9), .w(weight_reg22[15:8]), .out(acc_wire2_9), .resetn(resetn),.clk(clk));
PE PE2_10(.in(in_reg2_10), .acc(acc_reg1_10), .w(weight_reg22[23:16]), .out(acc_wire2_10), .resetn(resetn),.clk(clk));
PE PE2_11(.in(in_reg2_11), .acc(acc_reg1_11), .w(weight_reg22[31:24]), .out(acc_wire2_11), .resetn(resetn),.clk(clk));
PE PE2_12(.in(in_reg2_12), .acc(acc_reg1_12), .w(weight_reg23[7:0]), .out(acc_wire2_12), .resetn(resetn),.clk(clk));
PE PE2_13(.in(in_reg2_13), .acc(acc_reg1_13), .w(weight_reg23[15:8]), .out(acc_wire2_13), .resetn(resetn),.clk(clk));
PE PE2_14(.in(in_reg2_14), .acc(acc_reg1_14), .w(weight_reg23[23:16]), .out(acc_wire2_14), .resetn(resetn),.clk(clk));
PE PE2_15(.in(in_reg2_15), .acc(acc_reg1_15), .w(weight_reg23[31:24]), .out(acc_wire2_15), .resetn(resetn),.clk(clk));

PE PE3_0(.in(input3), .acc(acc_reg2_0), .w(weight_reg30[7:0]), .out(acc_wire3_0), .resetn(resetn),.clk(clk));
PE PE3_1(.in(in_reg3_1), .acc(acc_reg2_1), .w(weight_reg30[15:8]), .out(acc_wire3_1), .resetn(resetn),.clk(clk));
PE PE3_2(.in(in_reg3_2), .acc(acc_reg2_2), .w(weight_reg30[23:16]), .out(acc_wire3_2), .resetn(resetn),.clk(clk));
PE PE3_3(.in(in_reg3_3), .acc(acc_reg2_3), .w(weight_reg30[31:24]), .out(acc_wire3_3), .resetn(resetn),.clk(clk));
PE PE3_4(.in(in_reg3_4), .acc(acc_reg2_4), .w(weight_reg31[7:0]), .out(acc_wire3_4), .resetn(resetn),.clk(clk));
PE PE3_5(.in(in_reg3_5), .acc(acc_reg2_5), .w(weight_reg31[15:8]), .out(acc_wire3_5), .resetn(resetn),.clk(clk));
PE PE3_6(.in(in_reg3_6), .acc(acc_reg2_6), .w(weight_reg31[23:16]), .out(acc_wire3_6), .resetn(resetn),.clk(clk));
PE PE3_7(.in(in_reg3_7), .acc(acc_reg2_7), .w(weight_reg31[31:24]), .out(acc_wire3_7), .resetn(resetn),.clk(clk));
PE PE3_8(.in(in_reg3_8), .acc(acc_reg2_8), .w(weight_reg32[7:0]), .out(acc_wire3_8), .resetn(resetn),.clk(clk));
PE PE3_9(.in(in_reg3_9), .acc(acc_reg2_9), .w(weight_reg32[15:8]), .out(acc_wire3_9), .resetn(resetn),.clk(clk));
PE PE3_10(.in(in_reg3_10), .acc(acc_reg2_10), .w(weight_reg32[23:16]), .out(acc_wire3_10), .resetn(resetn),.clk(clk));
PE PE3_11(.in(in_reg3_11), .acc(acc_reg2_11), .w(weight_reg32[31:24]), .out(acc_wire3_11), .resetn(resetn),.clk(clk));
PE PE3_12(.in(in_reg3_12), .acc(acc_reg2_12), .w(weight_reg33[7:0]), .out(acc_wire3_12), .resetn(resetn),.clk(clk));
PE PE3_13(.in(in_reg3_13), .acc(acc_reg2_13), .w(weight_reg33[15:8]), .out(acc_wire3_13), .resetn(resetn),.clk(clk));
PE PE3_14(.in(in_reg3_14), .acc(acc_reg2_14), .w(weight_reg33[23:16]), .out(acc_wire3_14), .resetn(resetn),.clk(clk));
PE PE3_15(.in(in_reg3_15), .acc(acc_reg2_15), .w(weight_reg33[31:24]), .out(acc_wire3_15), .resetn(resetn),.clk(clk));

PE PE4_0(.in(input4), .acc(acc_reg3_0), .w(weight_reg40[7:0]), .out(acc_wire4_0), .resetn(resetn),.clk(clk));
PE PE4_1(.in(in_reg4_1), .acc(acc_reg3_1), .w(weight_reg40[15:8]), .out(acc_wire4_1), .resetn(resetn),.clk(clk));
PE PE4_2(.in(in_reg4_2), .acc(acc_reg3_2), .w(weight_reg40[23:16]), .out(acc_wire4_2), .resetn(resetn),.clk(clk));
PE PE4_3(.in(in_reg4_3), .acc(acc_reg3_3), .w(weight_reg40[31:24]), .out(acc_wire4_3), .resetn(resetn),.clk(clk));
PE PE4_4(.in(in_reg4_4), .acc(acc_reg3_4), .w(weight_reg41[7:0]), .out(acc_wire4_4), .resetn(resetn),.clk(clk));
PE PE4_5(.in(in_reg4_5), .acc(acc_reg3_5), .w(weight_reg41[15:8]), .out(acc_wire4_5), .resetn(resetn),.clk(clk));
PE PE4_6(.in(in_reg4_6), .acc(acc_reg3_6), .w(weight_reg41[23:16]), .out(acc_wire4_6), .resetn(resetn),.clk(clk));
PE PE4_7(.in(in_reg4_7), .acc(acc_reg3_7), .w(weight_reg41[31:24]), .out(acc_wire4_7), .resetn(resetn),.clk(clk));
PE PE4_8(.in(in_reg4_8), .acc(acc_reg3_8), .w(weight_reg42[7:0]), .out(acc_wire4_8), .resetn(resetn),.clk(clk));
PE PE4_9(.in(in_reg4_9), .acc(acc_reg3_9), .w(weight_reg42[15:8]), .out(acc_wire4_9), .resetn(resetn),.clk(clk));
PE PE4_10(.in(in_reg4_10), .acc(acc_reg3_10), .w(weight_reg42[23:16]), .out(acc_wire4_10), .resetn(resetn),.clk(clk));
PE PE4_11(.in(in_reg4_11), .acc(acc_reg3_11), .w(weight_reg42[31:24]), .out(acc_wire4_11), .resetn(resetn),.clk(clk));
PE PE4_12(.in(in_reg4_12), .acc(acc_reg3_12), .w(weight_reg43[7:0]), .out(acc_wire4_12), .resetn(resetn),.clk(clk));
PE PE4_13(.in(in_reg4_13), .acc(acc_reg3_13), .w(weight_reg43[15:8]), .out(acc_wire4_13), .resetn(resetn),.clk(clk));
PE PE4_14(.in(in_reg4_14), .acc(acc_reg3_14), .w(weight_reg43[23:16]), .out(acc_wire4_14), .resetn(resetn),.clk(clk));
PE PE4_15(.in(in_reg4_15), .acc(acc_reg3_15), .w(weight_reg43[31:24]), .out(acc_wire4_15), .resetn(resetn),.clk(clk));

PE PE5_0(.in(input5), .acc(acc_reg4_0), .w(weight_reg50[7:0]), .out(acc_wire5_0), .resetn(resetn),.clk(clk));
PE PE5_1(.in(in_reg5_1), .acc(acc_reg4_1), .w(weight_reg50[15:8]), .out(acc_wire5_1), .resetn(resetn),.clk(clk));
PE PE5_2(.in(in_reg5_2), .acc(acc_reg4_2), .w(weight_reg50[23:16]), .out(acc_wire5_2), .resetn(resetn),.clk(clk));
PE PE5_3(.in(in_reg5_3), .acc(acc_reg4_3), .w(weight_reg50[31:24]), .out(acc_wire5_3), .resetn(resetn),.clk(clk));
PE PE5_4(.in(in_reg5_4), .acc(acc_reg4_4), .w(weight_reg51[7:0]), .out(acc_wire5_4), .resetn(resetn),.clk(clk));
PE PE5_5(.in(in_reg5_5), .acc(acc_reg4_5), .w(weight_reg51[15:8]), .out(acc_wire5_5), .resetn(resetn),.clk(clk));
PE PE5_6(.in(in_reg5_6), .acc(acc_reg4_6), .w(weight_reg51[23:16]), .out(acc_wire5_6), .resetn(resetn),.clk(clk));
PE PE5_7(.in(in_reg5_7), .acc(acc_reg4_7), .w(weight_reg51[31:24]), .out(acc_wire5_7), .resetn(resetn),.clk(clk));
PE PE5_8(.in(in_reg5_8), .acc(acc_reg4_8), .w(weight_reg52[7:0]), .out(acc_wire5_8), .resetn(resetn),.clk(clk));
PE PE5_9(.in(in_reg5_9), .acc(acc_reg4_9), .w(weight_reg52[15:8]), .out(acc_wire5_9), .resetn(resetn),.clk(clk));
PE PE5_10(.in(in_reg5_10), .acc(acc_reg4_10), .w(weight_reg52[23:16]), .out(acc_wire5_10), .resetn(resetn),.clk(clk));
PE PE5_11(.in(in_reg5_11), .acc(acc_reg4_11), .w(weight_reg52[31:24]), .out(acc_wire5_11), .resetn(resetn),.clk(clk));
PE PE5_12(.in(in_reg5_12), .acc(acc_reg4_12), .w(weight_reg53[7:0]), .out(acc_wire5_12), .resetn(resetn),.clk(clk));
PE PE5_13(.in(in_reg5_13), .acc(acc_reg4_13), .w(weight_reg53[15:8]), .out(acc_wire5_13), .resetn(resetn),.clk(clk));
PE PE5_14(.in(in_reg5_14), .acc(acc_reg4_14), .w(weight_reg53[23:16]), .out(acc_wire5_14), .resetn(resetn),.clk(clk));
PE PE5_15(.in(in_reg5_15), .acc(acc_reg4_15), .w(weight_reg53[31:24]), .out(acc_wire5_15), .resetn(resetn),.clk(clk));

PE PE6_0(.in(input6), .acc(acc_reg5_0), .w(weight_reg60[7:0]), .out(acc_wire6_0), .resetn(resetn),.clk(clk));
PE PE6_1(.in(in_reg6_1), .acc(acc_reg5_1), .w(weight_reg60[15:8]), .out(acc_wire6_1), .resetn(resetn),.clk(clk));
PE PE6_2(.in(in_reg6_2), .acc(acc_reg5_2), .w(weight_reg60[23:16]), .out(acc_wire6_2), .resetn(resetn),.clk(clk));
PE PE6_3(.in(in_reg6_3), .acc(acc_reg5_3), .w(weight_reg60[31:24]), .out(acc_wire6_3), .resetn(resetn),.clk(clk));
PE PE6_4(.in(in_reg6_4), .acc(acc_reg5_4), .w(weight_reg61[7:0]), .out(acc_wire6_4), .resetn(resetn),.clk(clk));
PE PE6_5(.in(in_reg6_5), .acc(acc_reg5_5), .w(weight_reg61[15:8]), .out(acc_wire6_5), .resetn(resetn),.clk(clk));
PE PE6_6(.in(in_reg6_6), .acc(acc_reg5_6), .w(weight_reg61[23:16]), .out(acc_wire6_6), .resetn(resetn),.clk(clk));
PE PE6_7(.in(in_reg6_7), .acc(acc_reg5_7), .w(weight_reg61[31:24]), .out(acc_wire6_7), .resetn(resetn),.clk(clk));
PE PE6_8(.in(in_reg6_8), .acc(acc_reg5_8), .w(weight_reg62[7:0]), .out(acc_wire6_8), .resetn(resetn),.clk(clk));
PE PE6_9(.in(in_reg6_9), .acc(acc_reg5_9), .w(weight_reg62[15:8]), .out(acc_wire6_9), .resetn(resetn),.clk(clk));
PE PE6_10(.in(in_reg6_10), .acc(acc_reg5_10), .w(weight_reg62[23:16]), .out(acc_wire6_10), .resetn(resetn),.clk(clk));
PE PE6_11(.in(in_reg6_11), .acc(acc_reg5_11), .w(weight_reg62[31:24]), .out(acc_wire6_11), .resetn(resetn),.clk(clk));
PE PE6_12(.in(in_reg6_12), .acc(acc_reg5_12), .w(weight_reg63[7:0]), .out(acc_wire6_12), .resetn(resetn),.clk(clk));
PE PE6_13(.in(in_reg6_13), .acc(acc_reg5_13), .w(weight_reg63[15:8]), .out(acc_wire6_13), .resetn(resetn),.clk(clk));
PE PE6_14(.in(in_reg6_14), .acc(acc_reg5_14), .w(weight_reg63[23:16]), .out(acc_wire6_14), .resetn(resetn),.clk(clk));
PE PE6_15(.in(in_reg6_15), .acc(acc_reg5_15), .w(weight_reg63[31:24]), .out(acc_wire6_15), .resetn(resetn),.clk(clk));

PE PE7_0(.in(input7), .acc(acc_reg6_0), .w(weight_reg70[7:0]), .out(acc_wire7_0), .resetn(resetn),.clk(clk));
PE PE7_1(.in(in_reg7_1), .acc(acc_reg6_1), .w(weight_reg70[15:8]), .out(acc_wire7_1), .resetn(resetn),.clk(clk));
PE PE7_2(.in(in_reg7_2), .acc(acc_reg6_2), .w(weight_reg70[23:16]), .out(acc_wire7_2), .resetn(resetn),.clk(clk));
PE PE7_3(.in(in_reg7_3), .acc(acc_reg6_3), .w(weight_reg70[31:24]), .out(acc_wire7_3), .resetn(resetn),.clk(clk));
PE PE7_4(.in(in_reg7_4), .acc(acc_reg6_4), .w(weight_reg71[7:0]), .out(acc_wire7_4), .resetn(resetn),.clk(clk));
PE PE7_5(.in(in_reg7_5), .acc(acc_reg6_5), .w(weight_reg71[15:8]), .out(acc_wire7_5), .resetn(resetn),.clk(clk));
PE PE7_6(.in(in_reg7_6), .acc(acc_reg6_6), .w(weight_reg71[23:16]), .out(acc_wire7_6), .resetn(resetn),.clk(clk));
PE PE7_7(.in(in_reg7_7), .acc(acc_reg6_7), .w(weight_reg71[31:24]), .out(acc_wire7_7), .resetn(resetn),.clk(clk));
PE PE7_8(.in(in_reg7_8), .acc(acc_reg6_8), .w(weight_reg72[7:0]), .out(acc_wire7_8), .resetn(resetn),.clk(clk));
PE PE7_9(.in(in_reg7_9), .acc(acc_reg6_9), .w(weight_reg72[15:8]), .out(acc_wire7_9), .resetn(resetn),.clk(clk));
PE PE7_10(.in(in_reg7_10), .acc(acc_reg6_10), .w(weight_reg72[23:16]), .out(acc_wire7_10), .resetn(resetn),.clk(clk));
PE PE7_11(.in(in_reg7_11), .acc(acc_reg6_11), .w(weight_reg72[31:24]), .out(acc_wire7_11), .resetn(resetn),.clk(clk));
PE PE7_12(.in(in_reg7_12), .acc(acc_reg6_12), .w(weight_reg73[7:0]), .out(acc_wire7_12), .resetn(resetn),.clk(clk));
PE PE7_13(.in(in_reg7_13), .acc(acc_reg6_13), .w(weight_reg73[15:8]), .out(acc_wire7_13), .resetn(resetn),.clk(clk));
PE PE7_14(.in(in_reg7_14), .acc(acc_reg6_14), .w(weight_reg73[23:16]), .out(acc_wire7_14), .resetn(resetn),.clk(clk));
PE PE7_15(.in(in_reg7_15), .acc(acc_reg6_15), .w(weight_reg73[31:24]), .out(acc_wire7_15), .resetn(resetn),.clk(clk));

PE PE8_0(.in(input8), .acc(acc_reg7_0), .w(weight_reg80[7:0]), .out(acc_wire8_0), .resetn(resetn),.clk(clk));
PE PE8_1(.in(in_reg8_1), .acc(acc_reg7_1), .w(weight_reg80[15:8]), .out(acc_wire8_1), .resetn(resetn),.clk(clk));
PE PE8_2(.in(in_reg8_2), .acc(acc_reg7_2), .w(weight_reg80[23:16]), .out(acc_wire8_2), .resetn(resetn),.clk(clk));
PE PE8_3(.in(in_reg8_3), .acc(acc_reg7_3), .w(weight_reg80[31:24]), .out(acc_wire8_3), .resetn(resetn),.clk(clk));
PE PE8_4(.in(in_reg8_4), .acc(acc_reg7_4), .w(weight_reg81[7:0]), .out(acc_wire8_4), .resetn(resetn),.clk(clk));
PE PE8_5(.in(in_reg8_5), .acc(acc_reg7_5), .w(weight_reg81[15:8]), .out(acc_wire8_5), .resetn(resetn),.clk(clk));
PE PE8_6(.in(in_reg8_6), .acc(acc_reg7_6), .w(weight_reg81[23:16]), .out(acc_wire8_6), .resetn(resetn),.clk(clk));
PE PE8_7(.in(in_reg8_7), .acc(acc_reg7_7), .w(weight_reg81[31:24]), .out(acc_wire8_7), .resetn(resetn),.clk(clk));
PE PE8_8(.in(in_reg8_8), .acc(acc_reg7_8), .w(weight_reg82[7:0]), .out(acc_wire8_8), .resetn(resetn),.clk(clk));
PE PE8_9(.in(in_reg8_9), .acc(acc_reg7_9), .w(weight_reg82[15:8]), .out(acc_wire8_9), .resetn(resetn),.clk(clk));
PE PE8_10(.in(in_reg8_10), .acc(acc_reg7_10), .w(weight_reg82[23:16]), .out(acc_wire8_10), .resetn(resetn),.clk(clk));
PE PE8_11(.in(in_reg8_11), .acc(acc_reg7_11), .w(weight_reg82[31:24]), .out(acc_wire8_11), .resetn(resetn),.clk(clk));
PE PE8_12(.in(in_reg8_12), .acc(acc_reg7_12), .w(weight_reg83[7:0]), .out(acc_wire8_12), .resetn(resetn),.clk(clk));
PE PE8_13(.in(in_reg8_13), .acc(acc_reg7_13), .w(weight_reg83[15:8]), .out(acc_wire8_13), .resetn(resetn),.clk(clk));
PE PE8_14(.in(in_reg8_14), .acc(acc_reg7_14), .w(weight_reg83[23:16]), .out(acc_wire8_14), .resetn(resetn),.clk(clk));
PE PE8_15(.in(in_reg8_15), .acc(acc_reg7_15), .w(weight_reg83[31:24]), .out(acc_wire8_15), .resetn(resetn),.clk(clk));

PE PE9_0(.in(input9), .acc(acc_reg8_0), .w(weight_reg90[7:0]), .out(acc_wire9_0), .resetn(resetn),.clk(clk));
PE PE9_1(.in(in_reg9_1), .acc(acc_reg8_1), .w(weight_reg90[15:8]), .out(acc_wire9_1), .resetn(resetn),.clk(clk));
PE PE9_2(.in(in_reg9_2), .acc(acc_reg8_2), .w(weight_reg90[23:16]), .out(acc_wire9_2), .resetn(resetn),.clk(clk));
PE PE9_3(.in(in_reg9_3), .acc(acc_reg8_3), .w(weight_reg90[31:24]), .out(acc_wire9_3), .resetn(resetn),.clk(clk));
PE PE9_4(.in(in_reg9_4), .acc(acc_reg8_4), .w(weight_reg91[7:0]), .out(acc_wire9_4), .resetn(resetn),.clk(clk));
PE PE9_5(.in(in_reg9_5), .acc(acc_reg8_5), .w(weight_reg91[15:8]), .out(acc_wire9_5), .resetn(resetn),.clk(clk));
PE PE9_6(.in(in_reg9_6), .acc(acc_reg8_6), .w(weight_reg91[23:16]), .out(acc_wire9_6), .resetn(resetn),.clk(clk));
PE PE9_7(.in(in_reg9_7), .acc(acc_reg8_7), .w(weight_reg91[31:24]), .out(acc_wire9_7), .resetn(resetn),.clk(clk));
PE PE9_8(.in(in_reg9_8), .acc(acc_reg8_8), .w(weight_reg92[7:0]), .out(acc_wire9_8), .resetn(resetn),.clk(clk));
PE PE9_9(.in(in_reg9_9), .acc(acc_reg8_9), .w(weight_reg92[15:8]), .out(acc_wire9_9), .resetn(resetn),.clk(clk));
PE PE9_10(.in(in_reg9_10), .acc(acc_reg8_10), .w(weight_reg92[23:16]), .out(acc_wire9_10), .resetn(resetn),.clk(clk));
PE PE9_11(.in(in_reg9_11), .acc(acc_reg8_11), .w(weight_reg92[31:24]), .out(acc_wire9_11), .resetn(resetn),.clk(clk));
PE PE9_12(.in(in_reg9_12), .acc(acc_reg8_12), .w(weight_reg93[7:0]), .out(acc_wire9_12), .resetn(resetn),.clk(clk));
PE PE9_13(.in(in_reg9_13), .acc(acc_reg8_13), .w(weight_reg93[15:8]), .out(acc_wire9_13), .resetn(resetn),.clk(clk));
PE PE9_14(.in(in_reg9_14), .acc(acc_reg8_14), .w(weight_reg93[23:16]), .out(acc_wire9_14), .resetn(resetn),.clk(clk));
PE PE9_15(.in(in_reg9_15), .acc(acc_reg8_15), .w(weight_reg93[31:24]), .out(acc_wire9_15), .resetn(resetn),.clk(clk));

PE PE10_0(.in(input10), .acc(acc_reg9_0), .w(weight_reg100[7:0]), .out(acc_wire10_0), .resetn(resetn),.clk(clk));
PE PE10_1(.in(in_reg10_1), .acc(acc_reg9_1), .w(weight_reg100[15:8]), .out(acc_wire10_1), .resetn(resetn),.clk(clk));
PE PE10_2(.in(in_reg10_2), .acc(acc_reg9_2), .w(weight_reg100[23:16]), .out(acc_wire10_2), .resetn(resetn),.clk(clk));
PE PE10_3(.in(in_reg10_3), .acc(acc_reg9_3), .w(weight_reg100[31:24]), .out(acc_wire10_3), .resetn(resetn),.clk(clk));
PE PE10_4(.in(in_reg10_4), .acc(acc_reg9_4), .w(weight_reg101[7:0]), .out(acc_wire10_4), .resetn(resetn),.clk(clk));
PE PE10_5(.in(in_reg10_5), .acc(acc_reg9_5), .w(weight_reg101[15:8]), .out(acc_wire10_5), .resetn(resetn),.clk(clk));
PE PE10_6(.in(in_reg10_6), .acc(acc_reg9_6), .w(weight_reg101[23:16]), .out(acc_wire10_6), .resetn(resetn),.clk(clk));
PE PE10_7(.in(in_reg10_7), .acc(acc_reg9_7), .w(weight_reg101[31:24]), .out(acc_wire10_7), .resetn(resetn),.clk(clk));
PE PE10_8(.in(in_reg10_8), .acc(acc_reg9_8), .w(weight_reg102[7:0]), .out(acc_wire10_8), .resetn(resetn),.clk(clk));
PE PE10_9(.in(in_reg10_9), .acc(acc_reg9_9), .w(weight_reg102[15:8]), .out(acc_wire10_9), .resetn(resetn),.clk(clk));
PE PE10_10(.in(in_reg10_10), .acc(acc_reg9_10), .w(weight_reg102[23:16]), .out(acc_wire10_10), .resetn(resetn),.clk(clk));
PE PE10_11(.in(in_reg10_11), .acc(acc_reg9_11), .w(weight_reg102[31:24]), .out(acc_wire10_11), .resetn(resetn),.clk(clk));
PE PE10_12(.in(in_reg10_12), .acc(acc_reg9_12), .w(weight_reg103[7:0]), .out(acc_wire10_12), .resetn(resetn),.clk(clk));
PE PE10_13(.in(in_reg10_13), .acc(acc_reg9_13), .w(weight_reg103[15:8]), .out(acc_wire10_13), .resetn(resetn),.clk(clk));
PE PE10_14(.in(in_reg10_14), .acc(acc_reg9_14), .w(weight_reg103[23:16]), .out(acc_wire10_14), .resetn(resetn),.clk(clk));
PE PE10_15(.in(in_reg10_15), .acc(acc_reg9_15), .w(weight_reg103[31:24]), .out(acc_wire10_15), .resetn(resetn),.clk(clk));

PE PE11_0(.in(input11), .acc(acc_reg10_0), .w(weight_reg110[7:0]), .out(acc_wire11_0), .resetn(resetn),.clk(clk));
PE PE11_1(.in(in_reg11_1), .acc(acc_reg10_1), .w(weight_reg110[15:8]), .out(acc_wire11_1), .resetn(resetn),.clk(clk));
PE PE11_2(.in(in_reg11_2), .acc(acc_reg10_2), .w(weight_reg110[23:16]), .out(acc_wire11_2), .resetn(resetn),.clk(clk));
PE PE11_3(.in(in_reg11_3), .acc(acc_reg10_3), .w(weight_reg110[31:24]), .out(acc_wire11_3), .resetn(resetn),.clk(clk));
PE PE11_4(.in(in_reg11_4), .acc(acc_reg10_4), .w(weight_reg111[7:0]), .out(acc_wire11_4), .resetn(resetn),.clk(clk));
PE PE11_5(.in(in_reg11_5), .acc(acc_reg10_5), .w(weight_reg111[15:8]), .out(acc_wire11_5), .resetn(resetn),.clk(clk));
PE PE11_6(.in(in_reg11_6), .acc(acc_reg10_6), .w(weight_reg111[23:16]), .out(acc_wire11_6), .resetn(resetn),.clk(clk));
PE PE11_7(.in(in_reg11_7), .acc(acc_reg10_7), .w(weight_reg111[31:24]), .out(acc_wire11_7), .resetn(resetn),.clk(clk));
PE PE11_8(.in(in_reg11_8), .acc(acc_reg10_8), .w(weight_reg112[7:0]), .out(acc_wire11_8), .resetn(resetn),.clk(clk));
PE PE11_9(.in(in_reg11_9), .acc(acc_reg10_9), .w(weight_reg112[15:8]), .out(acc_wire11_9), .resetn(resetn),.clk(clk));
PE PE11_10(.in(in_reg11_10), .acc(acc_reg10_10), .w(weight_reg112[23:16]), .out(acc_wire11_10), .resetn(resetn),.clk(clk));
PE PE11_11(.in(in_reg11_11), .acc(acc_reg10_11), .w(weight_reg112[31:24]), .out(acc_wire11_11), .resetn(resetn),.clk(clk));
PE PE11_12(.in(in_reg11_12), .acc(acc_reg10_12), .w(weight_reg113[7:0]), .out(acc_wire11_12), .resetn(resetn),.clk(clk));
PE PE11_13(.in(in_reg11_13), .acc(acc_reg10_13), .w(weight_reg113[15:8]), .out(acc_wire11_13), .resetn(resetn),.clk(clk));
PE PE11_14(.in(in_reg11_14), .acc(acc_reg10_14), .w(weight_reg113[23:16]), .out(acc_wire11_14), .resetn(resetn),.clk(clk));
PE PE11_15(.in(in_reg11_15), .acc(acc_reg10_15), .w(weight_reg113[31:24]), .out(acc_wire11_15), .resetn(resetn),.clk(clk));

PE PE12_0(.in(input12), .acc(acc_reg11_0), .w(weight_reg120[7:0]), .out(acc_wire12_0), .resetn(resetn),.clk(clk));
PE PE12_1(.in(in_reg12_1), .acc(acc_reg11_1), .w(weight_reg120[15:8]), .out(acc_wire12_1), .resetn(resetn),.clk(clk));
PE PE12_2(.in(in_reg12_2), .acc(acc_reg11_2), .w(weight_reg120[23:16]), .out(acc_wire12_2), .resetn(resetn),.clk(clk));
PE PE12_3(.in(in_reg12_3), .acc(acc_reg11_3), .w(weight_reg120[31:24]), .out(acc_wire12_3), .resetn(resetn),.clk(clk));
PE PE12_4(.in(in_reg12_4), .acc(acc_reg11_4), .w(weight_reg121[7:0]), .out(acc_wire12_4), .resetn(resetn),.clk(clk));
PE PE12_5(.in(in_reg12_5), .acc(acc_reg11_5), .w(weight_reg121[15:8]), .out(acc_wire12_5), .resetn(resetn),.clk(clk));
PE PE12_6(.in(in_reg12_6), .acc(acc_reg11_6), .w(weight_reg121[23:16]), .out(acc_wire12_6), .resetn(resetn),.clk(clk));
PE PE12_7(.in(in_reg12_7), .acc(acc_reg11_7), .w(weight_reg121[31:24]), .out(acc_wire12_7), .resetn(resetn),.clk(clk));
PE PE12_8(.in(in_reg12_8), .acc(acc_reg11_8), .w(weight_reg122[7:0]), .out(acc_wire12_8), .resetn(resetn),.clk(clk));
PE PE12_9(.in(in_reg12_9), .acc(acc_reg11_9), .w(weight_reg122[15:8]), .out(acc_wire12_9), .resetn(resetn),.clk(clk));
PE PE12_10(.in(in_reg12_10), .acc(acc_reg11_10), .w(weight_reg122[23:16]), .out(acc_wire12_10), .resetn(resetn),.clk(clk));
PE PE12_11(.in(in_reg12_11), .acc(acc_reg11_11), .w(weight_reg122[31:24]), .out(acc_wire12_11), .resetn(resetn),.clk(clk));
PE PE12_12(.in(in_reg12_12), .acc(acc_reg11_12), .w(weight_reg123[7:0]), .out(acc_wire12_12), .resetn(resetn),.clk(clk));
PE PE12_13(.in(in_reg12_13), .acc(acc_reg11_13), .w(weight_reg123[15:8]), .out(acc_wire12_13), .resetn(resetn),.clk(clk));
PE PE12_14(.in(in_reg12_14), .acc(acc_reg11_14), .w(weight_reg123[23:16]), .out(acc_wire12_14), .resetn(resetn),.clk(clk));
PE PE12_15(.in(in_reg12_15), .acc(acc_reg11_15), .w(weight_reg123[31:24]), .out(acc_wire12_15), .resetn(resetn),.clk(clk));

PE PE13_0(.in(input13), .acc(acc_reg12_0), .w(weight_reg130[7:0]), .out(acc_wire13_0), .resetn(resetn),.clk(clk));
PE PE13_1(.in(in_reg13_1), .acc(acc_reg12_1), .w(weight_reg130[15:8]), .out(acc_wire13_1), .resetn(resetn),.clk(clk));
PE PE13_2(.in(in_reg13_2), .acc(acc_reg12_2), .w(weight_reg130[23:16]), .out(acc_wire13_2), .resetn(resetn),.clk(clk));
PE PE13_3(.in(in_reg13_3), .acc(acc_reg12_3), .w(weight_reg130[31:24]), .out(acc_wire13_3), .resetn(resetn),.clk(clk));
PE PE13_4(.in(in_reg13_4), .acc(acc_reg12_4), .w(weight_reg131[7:0]), .out(acc_wire13_4), .resetn(resetn),.clk(clk));
PE PE13_5(.in(in_reg13_5), .acc(acc_reg12_5), .w(weight_reg131[15:8]), .out(acc_wire13_5), .resetn(resetn),.clk(clk));
PE PE13_6(.in(in_reg13_6), .acc(acc_reg12_6), .w(weight_reg131[23:16]), .out(acc_wire13_6), .resetn(resetn),.clk(clk));
PE PE13_7(.in(in_reg13_7), .acc(acc_reg12_7), .w(weight_reg131[31:24]), .out(acc_wire13_7), .resetn(resetn),.clk(clk));
PE PE13_8(.in(in_reg13_8), .acc(acc_reg12_8), .w(weight_reg132[7:0]), .out(acc_wire13_8), .resetn(resetn),.clk(clk));
PE PE13_9(.in(in_reg13_9), .acc(acc_reg12_9), .w(weight_reg132[15:8]), .out(acc_wire13_9), .resetn(resetn),.clk(clk));
PE PE13_10(.in(in_reg13_10), .acc(acc_reg12_10), .w(weight_reg132[23:16]), .out(acc_wire13_10), .resetn(resetn),.clk(clk));
PE PE13_11(.in(in_reg13_11), .acc(acc_reg12_11), .w(weight_reg132[31:24]), .out(acc_wire13_11), .resetn(resetn),.clk(clk));
PE PE13_12(.in(in_reg13_12), .acc(acc_reg12_12), .w(weight_reg133[7:0]), .out(acc_wire13_12), .resetn(resetn),.clk(clk));
PE PE13_13(.in(in_reg13_13), .acc(acc_reg12_13), .w(weight_reg133[15:8]), .out(acc_wire13_13), .resetn(resetn),.clk(clk));
PE PE13_14(.in(in_reg13_14), .acc(acc_reg12_14), .w(weight_reg133[23:16]), .out(acc_wire13_14), .resetn(resetn),.clk(clk));
PE PE13_15(.in(in_reg13_15), .acc(acc_reg12_15), .w(weight_reg133[31:24]), .out(acc_wire13_15), .resetn(resetn),.clk(clk));

PE PE14_0(.in(input14), .acc(acc_reg13_0), .w(weight_reg140[7:0]), .out(acc_wire14_0), .resetn(resetn),.clk(clk));
PE PE14_1(.in(in_reg14_1), .acc(acc_reg13_1), .w(weight_reg140[15:8]), .out(acc_wire14_1), .resetn(resetn),.clk(clk));
PE PE14_2(.in(in_reg14_2), .acc(acc_reg13_2), .w(weight_reg140[23:16]), .out(acc_wire14_2), .resetn(resetn),.clk(clk));
PE PE14_3(.in(in_reg14_3), .acc(acc_reg13_3), .w(weight_reg140[31:24]), .out(acc_wire14_3), .resetn(resetn),.clk(clk));
PE PE14_4(.in(in_reg14_4), .acc(acc_reg13_4), .w(weight_reg141[7:0]), .out(acc_wire14_4), .resetn(resetn),.clk(clk));
PE PE14_5(.in(in_reg14_5), .acc(acc_reg13_5), .w(weight_reg141[15:8]), .out(acc_wire14_5), .resetn(resetn),.clk(clk));
PE PE14_6(.in(in_reg14_6), .acc(acc_reg13_6), .w(weight_reg141[23:16]), .out(acc_wire14_6), .resetn(resetn),.clk(clk));
PE PE14_7(.in(in_reg14_7), .acc(acc_reg13_7), .w(weight_reg141[31:24]), .out(acc_wire14_7), .resetn(resetn),.clk(clk));
PE PE14_8(.in(in_reg14_8), .acc(acc_reg13_8), .w(weight_reg142[7:0]), .out(acc_wire14_8), .resetn(resetn),.clk(clk));
PE PE14_9(.in(in_reg14_9), .acc(acc_reg13_9), .w(weight_reg142[15:8]), .out(acc_wire14_9), .resetn(resetn),.clk(clk));
PE PE14_10(.in(in_reg14_10), .acc(acc_reg13_10), .w(weight_reg142[23:16]), .out(acc_wire14_10), .resetn(resetn),.clk(clk));
PE PE14_11(.in(in_reg14_11), .acc(acc_reg13_11), .w(weight_reg142[31:24]), .out(acc_wire14_11), .resetn(resetn),.clk(clk));
PE PE14_12(.in(in_reg14_12), .acc(acc_reg13_12), .w(weight_reg143[7:0]), .out(acc_wire14_12), .resetn(resetn),.clk(clk));
PE PE14_13(.in(in_reg14_13), .acc(acc_reg13_13), .w(weight_reg143[15:8]), .out(acc_wire14_13), .resetn(resetn),.clk(clk));
PE PE14_14(.in(in_reg14_14), .acc(acc_reg13_14), .w(weight_reg143[23:16]), .out(acc_wire14_14), .resetn(resetn),.clk(clk));
PE PE14_15(.in(in_reg14_15), .acc(acc_reg13_15), .w(weight_reg143[31:24]), .out(acc_wire14_15), .resetn(resetn),.clk(clk));

PE PE15_0(.in(input15), .acc(acc_reg14_0), .w(weight_reg150[7:0]), .out(acc_wire15_0), .resetn(resetn),.clk(clk));
PE PE15_1(.in(in_reg15_1), .acc(acc_reg14_1), .w(weight_reg150[15:8]), .out(acc_wire15_1), .resetn(resetn),.clk(clk));
PE PE15_2(.in(in_reg15_2), .acc(acc_reg14_2), .w(weight_reg150[23:16]), .out(acc_wire15_2), .resetn(resetn),.clk(clk));
PE PE15_3(.in(in_reg15_3), .acc(acc_reg14_3), .w(weight_reg150[31:24]), .out(acc_wire15_3), .resetn(resetn),.clk(clk));
PE PE15_4(.in(in_reg15_4), .acc(acc_reg14_4), .w(weight_reg151[7:0]), .out(acc_wire15_4), .resetn(resetn),.clk(clk));
PE PE15_5(.in(in_reg15_5), .acc(acc_reg14_5), .w(weight_reg151[15:8]), .out(acc_wire15_5), .resetn(resetn),.clk(clk));
PE PE15_6(.in(in_reg15_6), .acc(acc_reg14_6), .w(weight_reg151[23:16]), .out(acc_wire15_6), .resetn(resetn),.clk(clk));
PE PE15_7(.in(in_reg15_7), .acc(acc_reg14_7), .w(weight_reg151[31:24]), .out(acc_wire15_7), .resetn(resetn),.clk(clk));
PE PE15_8(.in(in_reg15_8), .acc(acc_reg14_8), .w(weight_reg152[7:0]), .out(acc_wire15_8), .resetn(resetn),.clk(clk));
PE PE15_9(.in(in_reg15_9), .acc(acc_reg14_9), .w(weight_reg152[15:8]), .out(acc_wire15_9), .resetn(resetn),.clk(clk));
PE PE15_10(.in(in_reg15_10), .acc(acc_reg14_10), .w(weight_reg152[23:16]), .out(acc_wire15_10), .resetn(resetn),.clk(clk));
PE PE15_11(.in(in_reg15_11), .acc(acc_reg14_11), .w(weight_reg152[31:24]), .out(acc_wire15_11), .resetn(resetn),.clk(clk));
PE PE15_12(.in(in_reg15_12), .acc(acc_reg14_12), .w(weight_reg153[7:0]), .out(acc_wire15_12), .resetn(resetn),.clk(clk));
PE PE15_13(.in(in_reg15_13), .acc(acc_reg14_13), .w(weight_reg153[15:8]), .out(acc_wire15_13), .resetn(resetn),.clk(clk));
PE PE15_14(.in(in_reg15_14), .acc(acc_reg14_14), .w(weight_reg153[23:16]), .out(acc_wire15_14), .resetn(resetn),.clk(clk));
PE PE15_15(.in(in_reg15_15), .acc(acc_reg14_15), .w(weight_reg153[31:24]), .out(acc_wire15_15), .resetn(resetn),.clk(clk));

wire calc_enable;
assign calc_enable = (col ==2'b11) && (command == 2'b10);
always@ (posedge clk)
begin
	if (calc_enable)
	begin
		in_reg0_1<= input0;
		in_reg1_1<= input1;
		in_reg2_1<= input2;
		in_reg3_1<= input3;
		in_reg4_1<= input4;
		in_reg5_1<= input5;
		in_reg6_1<= input6;
		in_reg7_1<= input7;
		in_reg8_1<= input8;
		in_reg9_1<= input9;
		in_reg10_1<= input10;
		in_reg11_1<= input11;
		in_reg12_1<= input12;
		in_reg13_1<= input13;
		in_reg14_1<= input14;
		in_reg15_1<= input15;
		
		in_reg0_2<= in_reg0_1;
		in_reg0_3<= in_reg0_2;
		in_reg0_4<= in_reg0_3;
		in_reg0_5<= in_reg0_4;
		in_reg0_6<= in_reg0_5;
		in_reg0_7<= in_reg0_6;
		in_reg0_8<= in_reg0_7;
		in_reg0_9<= in_reg0_8;
		in_reg0_10<= in_reg0_9;
		in_reg0_11<= in_reg0_10;
		in_reg0_12<= in_reg0_11;
		in_reg0_13<= in_reg0_12;
		in_reg0_14<= in_reg0_13;
		in_reg0_15<= in_reg0_14;
		in_reg1_2<= in_reg1_1;
		in_reg1_3<= in_reg1_2;
		in_reg1_4<= in_reg1_3;
		in_reg1_5<= in_reg1_4;
		in_reg1_6<= in_reg1_5;
		in_reg1_7<= in_reg1_6;
		in_reg1_8<= in_reg1_7;
		in_reg1_9<= in_reg1_8;
		in_reg1_10<= in_reg1_9;
		in_reg1_11<= in_reg1_10;
		in_reg1_12<= in_reg1_11;
		in_reg1_13<= in_reg1_12;
		in_reg1_14<= in_reg1_13;
		in_reg1_15<= in_reg1_14;
		in_reg2_2<= in_reg2_1;
		in_reg2_3<= in_reg2_2;
		in_reg2_4<= in_reg2_3;
		in_reg2_5<= in_reg2_4;
		in_reg2_6<= in_reg2_5;
		in_reg2_7<= in_reg2_6;
		in_reg2_8<= in_reg2_7;
		in_reg2_9<= in_reg2_8;
		in_reg2_10<= in_reg2_9;
		in_reg2_11<= in_reg2_10;
		in_reg2_12<= in_reg2_11;
		in_reg2_13<= in_reg2_12;
		in_reg2_14<= in_reg2_13;
		in_reg2_15<= in_reg2_14;
		in_reg3_2<= in_reg3_1;
		in_reg3_3<= in_reg3_2;
		in_reg3_4<= in_reg3_3;
		in_reg3_5<= in_reg3_4;
		in_reg3_6<= in_reg3_5;
		in_reg3_7<= in_reg3_6;
		in_reg3_8<= in_reg3_7;
		in_reg3_9<= in_reg3_8;
		in_reg3_10<= in_reg3_9;
		in_reg3_11<= in_reg3_10;
		in_reg3_12<= in_reg3_11;
		in_reg3_13<= in_reg3_12;
		in_reg3_14<= in_reg3_13;
		in_reg3_15<= in_reg3_14;
		in_reg4_2<= in_reg4_1;
		in_reg4_3<= in_reg4_2;
		in_reg4_4<= in_reg4_3;
		in_reg4_5<= in_reg4_4;
		in_reg4_6<= in_reg4_5;
		in_reg4_7<= in_reg4_6;
		in_reg4_8<= in_reg4_7;
		in_reg4_9<= in_reg4_8;
		in_reg4_10<= in_reg4_9;
		in_reg4_11<= in_reg4_10;
		in_reg4_12<= in_reg4_11;
		in_reg4_13<= in_reg4_12;
		in_reg4_14<= in_reg4_13;
		in_reg4_15<= in_reg4_14;
		in_reg5_2<= in_reg5_1;
		in_reg5_3<= in_reg5_2;
		in_reg5_4<= in_reg5_3;
		in_reg5_5<= in_reg5_4;
		in_reg5_6<= in_reg5_5;
		in_reg5_7<= in_reg5_6;
		in_reg5_8<= in_reg5_7;
		in_reg5_9<= in_reg5_8;
		in_reg5_10<= in_reg5_9;
		in_reg5_11<= in_reg5_10;
		in_reg5_12<= in_reg5_11;
		in_reg5_13<= in_reg5_12;
		in_reg5_14<= in_reg5_13;
		in_reg5_15<= in_reg5_14;
		in_reg6_2<= in_reg6_1;
		in_reg6_3<= in_reg6_2;
		in_reg6_4<= in_reg6_3;
		in_reg6_5<= in_reg6_4;
		in_reg6_6<= in_reg6_5;
		in_reg6_7<= in_reg6_6;
		in_reg6_8<= in_reg6_7;
		in_reg6_9<= in_reg6_8;
		in_reg6_10<= in_reg6_9;
		in_reg6_11<= in_reg6_10;
		in_reg6_12<= in_reg6_11;
		in_reg6_13<= in_reg6_12;
		in_reg6_14<= in_reg6_13;
		in_reg6_15<= in_reg6_14;
		in_reg7_2<= in_reg7_1;
		in_reg7_3<= in_reg7_2;
		in_reg7_4<= in_reg7_3;
		in_reg7_5<= in_reg7_4;
		in_reg7_6<= in_reg7_5;
		in_reg7_7<= in_reg7_6;
		in_reg7_8<= in_reg7_7;
		in_reg7_9<= in_reg7_8;
		in_reg7_10<= in_reg7_9;
		in_reg7_11<= in_reg7_10;
		in_reg7_12<= in_reg7_11;
		in_reg7_13<= in_reg7_12;
		in_reg7_14<= in_reg7_13;
		in_reg7_15<= in_reg7_14;
		in_reg8_2<= in_reg8_1;
		in_reg8_3<= in_reg8_2;
		in_reg8_4<= in_reg8_3;
		in_reg8_5<= in_reg8_4;
		in_reg8_6<= in_reg8_5;
		in_reg8_7<= in_reg8_6;
		in_reg8_8<= in_reg8_7;
		in_reg8_9<= in_reg8_8;
		in_reg8_10<= in_reg8_9;
		in_reg8_11<= in_reg8_10;
		in_reg8_12<= in_reg8_11;
		in_reg8_13<= in_reg8_12;
		in_reg8_14<= in_reg8_13;
		in_reg8_15<= in_reg8_14;
		in_reg9_2<= in_reg9_1;
		in_reg9_3<= in_reg9_2;
		in_reg9_4<= in_reg9_3;
		in_reg9_5<= in_reg9_4;
		in_reg9_6<= in_reg9_5;
		in_reg9_7<= in_reg9_6;
		in_reg9_8<= in_reg9_7;
		in_reg9_9<= in_reg9_8;
		in_reg9_10<= in_reg9_9;
		in_reg9_11<= in_reg9_10;
		in_reg9_12<= in_reg9_11;
		in_reg9_13<= in_reg9_12;
		in_reg9_14<= in_reg9_13;
		in_reg9_15<= in_reg9_14;
		in_reg10_2<= in_reg10_1;
		in_reg10_3<= in_reg10_2;
		in_reg10_4<= in_reg10_3;
		in_reg10_5<= in_reg10_4;
		in_reg10_6<= in_reg10_5;
		in_reg10_7<= in_reg10_6;
		in_reg10_8<= in_reg10_7;
		in_reg10_9<= in_reg10_8;
		in_reg10_10<= in_reg10_9;
		in_reg10_11<= in_reg10_10;
		in_reg10_12<= in_reg10_11;
		in_reg10_13<= in_reg10_12;
		in_reg10_14<= in_reg10_13;
		in_reg10_15<= in_reg10_14;
		in_reg11_2<= in_reg11_1;
		in_reg11_3<= in_reg11_2;
		in_reg11_4<= in_reg11_3;
		in_reg11_5<= in_reg11_4;
		in_reg11_6<= in_reg11_5;
		in_reg11_7<= in_reg11_6;
		in_reg11_8<= in_reg11_7;
		in_reg11_9<= in_reg11_8;
		in_reg11_10<= in_reg11_9;
		in_reg11_11<= in_reg11_10;
		in_reg11_12<= in_reg11_11;
		in_reg11_13<= in_reg11_12;
		in_reg11_14<= in_reg11_13;
		in_reg11_15<= in_reg11_14;
		in_reg12_2<= in_reg12_1;
		in_reg12_3<= in_reg12_2;
		in_reg12_4<= in_reg12_3;
		in_reg12_5<= in_reg12_4;
		in_reg12_6<= in_reg12_5;
		in_reg12_7<= in_reg12_6;
		in_reg12_8<= in_reg12_7;
		in_reg12_9<= in_reg12_8;
		in_reg12_10<= in_reg12_9;
		in_reg12_11<= in_reg12_10;
		in_reg12_12<= in_reg12_11;
		in_reg12_13<= in_reg12_12;
		in_reg12_14<= in_reg12_13;
		in_reg12_15<= in_reg12_14;
		in_reg13_2<= in_reg13_1;
		in_reg13_3<= in_reg13_2;
		in_reg13_4<= in_reg13_3;
		in_reg13_5<= in_reg13_4;
		in_reg13_6<= in_reg13_5;
		in_reg13_7<= in_reg13_6;
		in_reg13_8<= in_reg13_7;
		in_reg13_9<= in_reg13_8;
		in_reg13_10<= in_reg13_9;
		in_reg13_11<= in_reg13_10;
		in_reg13_12<= in_reg13_11;
		in_reg13_13<= in_reg13_12;
		in_reg13_14<= in_reg13_13;
		in_reg13_15<= in_reg13_14;
		in_reg14_2<= in_reg14_1;
		in_reg14_3<= in_reg14_2;
		in_reg14_4<= in_reg14_3;
		in_reg14_5<= in_reg14_4;
		in_reg14_6<= in_reg14_5;
		in_reg14_7<= in_reg14_6;
		in_reg14_8<= in_reg14_7;
		in_reg14_9<= in_reg14_8;
		in_reg14_10<= in_reg14_9;
		in_reg14_11<= in_reg14_10;
		in_reg14_12<= in_reg14_11;
		in_reg14_13<= in_reg14_12;
		in_reg14_14<= in_reg14_13;
		in_reg14_15<= in_reg14_14;
		in_reg15_2<= in_reg15_1;
		in_reg15_3<= in_reg15_2;
		in_reg15_4<= in_reg15_3;
		in_reg15_5<= in_reg15_4;
		in_reg15_6<= in_reg15_5;
		in_reg15_7<= in_reg15_6;
		in_reg15_8<= in_reg15_7;
		in_reg15_9<= in_reg15_8;
		in_reg15_10<= in_reg15_9;
		in_reg15_11<= in_reg15_10;
		in_reg15_12<= in_reg15_11;
		in_reg15_13<= in_reg15_12;
		in_reg15_14<= in_reg15_13;
		in_reg15_15<= in_reg15_14;
	end
end

always@ (posedge clk)
begin
	if (calc_enable)
	begin
		acc_reg0_0 <= acc_wire0_0;
		acc_reg0_1 <= acc_wire0_1;
		acc_reg0_2 <= acc_wire0_2;
		acc_reg0_3 <= acc_wire0_3;
		acc_reg0_4 <= acc_wire0_4;
		acc_reg0_5 <= acc_wire0_5;
		acc_reg0_6 <= acc_wire0_6;
		acc_reg0_7 <= acc_wire0_7;
		acc_reg0_8 <= acc_wire0_8;
		acc_reg0_9 <= acc_wire0_9;
		acc_reg0_10 <= acc_wire0_10;
		acc_reg0_11 <= acc_wire0_11;
		acc_reg0_12 <= acc_wire0_12;
		acc_reg0_13 <= acc_wire0_13;
		acc_reg0_14 <= acc_wire0_14;
		acc_reg0_15 <= acc_wire0_15;
		acc_reg1_0 <= acc_wire1_0;
		acc_reg1_1 <= acc_wire1_1;
		acc_reg1_2 <= acc_wire1_2;
		acc_reg1_3 <= acc_wire1_3;
		acc_reg1_4 <= acc_wire1_4;
		acc_reg1_5 <= acc_wire1_5;
		acc_reg1_6 <= acc_wire1_6;
		acc_reg1_7 <= acc_wire1_7;
		acc_reg1_8 <= acc_wire1_8;
		acc_reg1_9 <= acc_wire1_9;
		acc_reg1_10 <= acc_wire1_10;
		acc_reg1_11 <= acc_wire1_11;
		acc_reg1_12 <= acc_wire1_12;
		acc_reg1_13 <= acc_wire1_13;
		acc_reg1_14 <= acc_wire1_14;
		acc_reg1_15 <= acc_wire1_15;
		acc_reg2_0 <= acc_wire2_0;
		acc_reg2_1 <= acc_wire2_1;
		acc_reg2_2 <= acc_wire2_2;
		acc_reg2_3 <= acc_wire2_3;
		acc_reg2_4 <= acc_wire2_4;
		acc_reg2_5 <= acc_wire2_5;
		acc_reg2_6 <= acc_wire2_6;
		acc_reg2_7 <= acc_wire2_7;
		acc_reg2_8 <= acc_wire2_8;
		acc_reg2_9 <= acc_wire2_9;
		acc_reg2_10 <= acc_wire2_10;
		acc_reg2_11 <= acc_wire2_11;
		acc_reg2_12 <= acc_wire2_12;
		acc_reg2_13 <= acc_wire2_13;
		acc_reg2_14 <= acc_wire2_14;
		acc_reg2_15 <= acc_wire2_15;
		acc_reg3_0 <= acc_wire3_0;
		acc_reg3_1 <= acc_wire3_1;
		acc_reg3_2 <= acc_wire3_2;
		acc_reg3_3 <= acc_wire3_3;
		acc_reg3_4 <= acc_wire3_4;
		acc_reg3_5 <= acc_wire3_5;
		acc_reg3_6 <= acc_wire3_6;
		acc_reg3_7 <= acc_wire3_7;
		acc_reg3_8 <= acc_wire3_8;
		acc_reg3_9 <= acc_wire3_9;
		acc_reg3_10 <= acc_wire3_10;
		acc_reg3_11 <= acc_wire3_11;
		acc_reg3_12 <= acc_wire3_12;
		acc_reg3_13 <= acc_wire3_13;
		acc_reg3_14 <= acc_wire3_14;
		acc_reg3_15 <= acc_wire3_15;
		acc_reg4_0 <= acc_wire4_0;
		acc_reg4_1 <= acc_wire4_1;
		acc_reg4_2 <= acc_wire4_2;
		acc_reg4_3 <= acc_wire4_3;
		acc_reg4_4 <= acc_wire4_4;
		acc_reg4_5 <= acc_wire4_5;
		acc_reg4_6 <= acc_wire4_6;
		acc_reg4_7 <= acc_wire4_7;
		acc_reg4_8 <= acc_wire4_8;
		acc_reg4_9 <= acc_wire4_9;
		acc_reg4_10 <= acc_wire4_10;
		acc_reg4_11 <= acc_wire4_11;
		acc_reg4_12 <= acc_wire4_12;
		acc_reg4_13 <= acc_wire4_13;
		acc_reg4_14 <= acc_wire4_14;
		acc_reg4_15 <= acc_wire4_15;
		acc_reg5_0 <= acc_wire5_0;
		acc_reg5_1 <= acc_wire5_1;
		acc_reg5_2 <= acc_wire5_2;
		acc_reg5_3 <= acc_wire5_3;
		acc_reg5_4 <= acc_wire5_4;
		acc_reg5_5 <= acc_wire5_5;
		acc_reg5_6 <= acc_wire5_6;
		acc_reg5_7 <= acc_wire5_7;
		acc_reg5_8 <= acc_wire5_8;
		acc_reg5_9 <= acc_wire5_9;
		acc_reg5_10 <= acc_wire5_10;
		acc_reg5_11 <= acc_wire5_11;
		acc_reg5_12 <= acc_wire5_12;
		acc_reg5_13 <= acc_wire5_13;
		acc_reg5_14 <= acc_wire5_14;
		acc_reg5_15 <= acc_wire5_15;
		acc_reg6_0 <= acc_wire6_0;
		acc_reg6_1 <= acc_wire6_1;
		acc_reg6_2 <= acc_wire6_2;
		acc_reg6_3 <= acc_wire6_3;
		acc_reg6_4 <= acc_wire6_4;
		acc_reg6_5 <= acc_wire6_5;
		acc_reg6_6 <= acc_wire6_6;
		acc_reg6_7 <= acc_wire6_7;
		acc_reg6_8 <= acc_wire6_8;
		acc_reg6_9 <= acc_wire6_9;
		acc_reg6_10 <= acc_wire6_10;
		acc_reg6_11 <= acc_wire6_11;
		acc_reg6_12 <= acc_wire6_12;
		acc_reg6_13 <= acc_wire6_13;
		acc_reg6_14 <= acc_wire6_14;
		acc_reg6_15 <= acc_wire6_15;
		acc_reg7_0 <= acc_wire7_0;
		acc_reg7_1 <= acc_wire7_1;
		acc_reg7_2 <= acc_wire7_2;
		acc_reg7_3 <= acc_wire7_3;
		acc_reg7_4 <= acc_wire7_4;
		acc_reg7_5 <= acc_wire7_5;
		acc_reg7_6 <= acc_wire7_6;
		acc_reg7_7 <= acc_wire7_7;
		acc_reg7_8 <= acc_wire7_8;
		acc_reg7_9 <= acc_wire7_9;
		acc_reg7_10 <= acc_wire7_10;
		acc_reg7_11 <= acc_wire7_11;
		acc_reg7_12 <= acc_wire7_12;
		acc_reg7_13 <= acc_wire7_13;
		acc_reg7_14 <= acc_wire7_14;
		acc_reg7_15 <= acc_wire7_15;
		acc_reg8_0 <= acc_wire8_0;
		acc_reg8_1 <= acc_wire8_1;
		acc_reg8_2 <= acc_wire8_2;
		acc_reg8_3 <= acc_wire8_3;
		acc_reg8_4 <= acc_wire8_4;
		acc_reg8_5 <= acc_wire8_5;
		acc_reg8_6 <= acc_wire8_6;
		acc_reg8_7 <= acc_wire8_7;
		acc_reg8_8 <= acc_wire8_8;
		acc_reg8_9 <= acc_wire8_9;
		acc_reg8_10 <= acc_wire8_10;
		acc_reg8_11 <= acc_wire8_11;
		acc_reg8_12 <= acc_wire8_12;
		acc_reg8_13 <= acc_wire8_13;
		acc_reg8_14 <= acc_wire8_14;
		acc_reg8_15 <= acc_wire8_15;
		acc_reg9_0 <= acc_wire9_0;
		acc_reg9_1 <= acc_wire9_1;
		acc_reg9_2 <= acc_wire9_2;
		acc_reg9_3 <= acc_wire9_3;
		acc_reg9_4 <= acc_wire9_4;
		acc_reg9_5 <= acc_wire9_5;
		acc_reg9_6 <= acc_wire9_6;
		acc_reg9_7 <= acc_wire9_7;
		acc_reg9_8 <= acc_wire9_8;
		acc_reg9_9 <= acc_wire9_9;
		acc_reg9_10 <= acc_wire9_10;
		acc_reg9_11 <= acc_wire9_11;
		acc_reg9_12 <= acc_wire9_12;
		acc_reg9_13 <= acc_wire9_13;
		acc_reg9_14 <= acc_wire9_14;
		acc_reg9_15 <= acc_wire9_15;
		acc_reg10_0 <= acc_wire10_0;
		acc_reg10_1 <= acc_wire10_1;
		acc_reg10_2 <= acc_wire10_2;
		acc_reg10_3 <= acc_wire10_3;
		acc_reg10_4 <= acc_wire10_4;
		acc_reg10_5 <= acc_wire10_5;
		acc_reg10_6 <= acc_wire10_6;
		acc_reg10_7 <= acc_wire10_7;
		acc_reg10_8 <= acc_wire10_8;
		acc_reg10_9 <= acc_wire10_9;
		acc_reg10_10 <= acc_wire10_10;
		acc_reg10_11 <= acc_wire10_11;
		acc_reg10_12 <= acc_wire10_12;
		acc_reg10_13 <= acc_wire10_13;
		acc_reg10_14 <= acc_wire10_14;
		acc_reg10_15 <= acc_wire10_15;
		acc_reg11_0 <= acc_wire11_0;
		acc_reg11_1 <= acc_wire11_1;
		acc_reg11_2 <= acc_wire11_2;
		acc_reg11_3 <= acc_wire11_3;
		acc_reg11_4 <= acc_wire11_4;
		acc_reg11_5 <= acc_wire11_5;
		acc_reg11_6 <= acc_wire11_6;
		acc_reg11_7 <= acc_wire11_7;
		acc_reg11_8 <= acc_wire11_8;
		acc_reg11_9 <= acc_wire11_9;
		acc_reg11_10 <= acc_wire11_10;
		acc_reg11_11 <= acc_wire11_11;
		acc_reg11_12 <= acc_wire11_12;
		acc_reg11_13 <= acc_wire11_13;
		acc_reg11_14 <= acc_wire11_14;
		acc_reg11_15 <= acc_wire11_15;
		acc_reg12_0 <= acc_wire12_0;
		acc_reg12_1 <= acc_wire12_1;
		acc_reg12_2 <= acc_wire12_2;
		acc_reg12_3 <= acc_wire12_3;
		acc_reg12_4 <= acc_wire12_4;
		acc_reg12_5 <= acc_wire12_5;
		acc_reg12_6 <= acc_wire12_6;
		acc_reg12_7 <= acc_wire12_7;
		acc_reg12_8 <= acc_wire12_8;
		acc_reg12_9 <= acc_wire12_9;
		acc_reg12_10 <= acc_wire12_10;
		acc_reg12_11 <= acc_wire12_11;
		acc_reg12_12 <= acc_wire12_12;
		acc_reg12_13 <= acc_wire12_13;
		acc_reg12_14 <= acc_wire12_14;
		acc_reg12_15 <= acc_wire12_15;
		acc_reg13_0 <= acc_wire13_0;
		acc_reg13_1 <= acc_wire13_1;
		acc_reg13_2 <= acc_wire13_2;
		acc_reg13_3 <= acc_wire13_3;
		acc_reg13_4 <= acc_wire13_4;
		acc_reg13_5 <= acc_wire13_5;
		acc_reg13_6 <= acc_wire13_6;
		acc_reg13_7 <= acc_wire13_7;
		acc_reg13_8 <= acc_wire13_8;
		acc_reg13_9 <= acc_wire13_9;
		acc_reg13_10 <= acc_wire13_10;
		acc_reg13_11 <= acc_wire13_11;
		acc_reg13_12 <= acc_wire13_12;
		acc_reg13_13 <= acc_wire13_13;
		acc_reg13_14 <= acc_wire13_14;
		acc_reg13_15 <= acc_wire13_15;
		acc_reg14_0 <= acc_wire14_0;
		acc_reg14_1 <= acc_wire14_1;
		acc_reg14_2 <= acc_wire14_2;
		acc_reg14_3 <= acc_wire14_3;
		acc_reg14_4 <= acc_wire14_4;
		acc_reg14_5 <= acc_wire14_5;
		acc_reg14_6 <= acc_wire14_6;
		acc_reg14_7 <= acc_wire14_7;
		acc_reg14_8 <= acc_wire14_8;
		acc_reg14_9 <= acc_wire14_9;
		acc_reg14_10 <= acc_wire14_10;
		acc_reg14_11 <= acc_wire14_11;
		acc_reg14_12 <= acc_wire14_12;
		acc_reg14_13 <= acc_wire14_13;
		acc_reg14_14 <= acc_wire14_14;
		acc_reg14_15 <= acc_wire14_15;
		acc_reg15_0 <= acc_wire15_0;
		acc_reg15_1 <= acc_wire15_1;
		acc_reg15_2 <= acc_wire15_2;
		acc_reg15_3 <= acc_wire15_3;
		acc_reg15_4 <= acc_wire15_4;
		acc_reg15_5 <= acc_wire15_5;
		acc_reg15_6 <= acc_wire15_6;
		acc_reg15_7 <= acc_wire15_7;
		acc_reg15_8 <= acc_wire15_8;
		acc_reg15_9 <= acc_wire15_9;
		acc_reg15_10 <= acc_wire15_10;
		acc_reg15_11 <= acc_wire15_11;
		acc_reg15_12 <= acc_wire15_12;
		acc_reg15_13 <= acc_wire15_13;
		acc_reg15_14 <= acc_wire15_14;
		acc_reg15_15 <= acc_wire15_15;
	end
end
	
assign output0 = acc_reg15_0;
assign output1 = acc_reg15_1;
assign output2 = acc_reg15_2;
assign output3 = acc_reg15_3;
assign output4 = acc_reg15_4;
assign output5 = acc_reg15_5;
assign output6 = acc_reg15_6;
assign output7 = acc_reg15_7;
assign output8 = acc_reg15_8;
assign output9 = acc_reg15_9;
assign output10 = acc_reg15_10;
assign output11 = acc_reg15_11;
assign output12 = acc_reg15_12;
assign output13 = acc_reg15_13;
assign output14 = acc_reg15_14;
assign output15 = acc_reg15_15;

endmodule 
